magic
tech sky130A
magscale 1 2
timestamp 1672339081
<< viali >>
rect 2145 27557 2179 27591
rect 2789 27557 2823 27591
rect 3985 27557 4019 27591
rect 4629 27557 4663 27591
rect 6009 27557 6043 27591
rect 7113 27557 7147 27591
rect 8585 27557 8619 27591
rect 9597 27557 9631 27591
rect 11161 27557 11195 27591
rect 12081 27557 12115 27591
rect 14289 27557 14323 27591
rect 14933 27557 14967 27591
rect 16865 27557 16899 27591
rect 17509 27557 17543 27591
rect 18705 27557 18739 27591
rect 19533 27557 19567 27591
rect 21189 27557 21223 27591
rect 22017 27557 22051 27591
rect 1593 26945 1627 26979
rect 2237 26945 2271 26979
rect 22293 26809 22327 26843
rect 1593 26333 1627 26367
rect 22293 26333 22327 26367
rect 1593 25653 1627 25687
rect 22293 25245 22327 25279
rect 22293 24633 22327 24667
rect 1593 24157 1627 24191
rect 22293 23545 22327 23579
rect 1593 23477 1627 23511
rect 22293 23069 22327 23103
rect 1593 22389 1627 22423
rect 22293 22117 22327 22151
rect 1593 21437 1627 21471
rect 22293 21369 22327 21403
rect 22293 20281 22327 20315
rect 1593 20213 1627 20247
rect 1593 19805 1627 19839
rect 22293 19805 22327 19839
rect 22293 18717 22327 18751
rect 22293 18105 22327 18139
rect 1593 18037 1627 18071
rect 1593 17629 1627 17663
rect 22293 17017 22327 17051
rect 22293 16609 22327 16643
rect 1593 15997 1627 16031
rect 1593 15453 1627 15487
rect 22293 15453 22327 15487
rect 22293 14841 22327 14875
rect 1593 14365 1627 14399
rect 22293 13821 22327 13855
rect 1593 13277 1627 13311
rect 22293 13277 22327 13311
rect 1593 12189 1627 12223
rect 22293 12189 22327 12223
rect 22293 11577 22327 11611
rect 1593 11509 1627 11543
rect 22293 10489 22327 10523
rect 1593 10013 1627 10047
rect 22293 10013 22327 10047
rect 1593 9333 1627 9367
rect 22293 8925 22327 8959
rect 22293 8313 22327 8347
rect 1593 7837 1627 7871
rect 22293 7225 22327 7259
rect 1593 7157 1627 7191
rect 22293 6749 22327 6783
rect 1593 6069 1627 6103
rect 22293 5661 22327 5695
rect 1593 5117 1627 5151
rect 22293 5049 22327 5083
rect 22293 3961 22327 3995
rect 1593 3893 1627 3927
rect 1593 3485 1627 3519
rect 22293 3485 22327 3519
rect 1593 2805 1627 2839
rect 1593 2397 1627 2431
<< metal1 >>
rect 1104 27770 22816 27792
rect 1104 27718 3664 27770
rect 3716 27718 3728 27770
rect 3780 27718 3792 27770
rect 3844 27718 3856 27770
rect 3908 27718 3920 27770
rect 3972 27718 9092 27770
rect 9144 27718 9156 27770
rect 9208 27718 9220 27770
rect 9272 27718 9284 27770
rect 9336 27718 9348 27770
rect 9400 27718 14520 27770
rect 14572 27718 14584 27770
rect 14636 27718 14648 27770
rect 14700 27718 14712 27770
rect 14764 27718 14776 27770
rect 14828 27718 19948 27770
rect 20000 27718 20012 27770
rect 20064 27718 20076 27770
rect 20128 27718 20140 27770
rect 20192 27718 20204 27770
rect 20256 27718 22816 27770
rect 1104 27696 22816 27718
rect 2130 27588 2136 27600
rect 2091 27560 2136 27588
rect 2130 27548 2136 27560
rect 2188 27548 2194 27600
rect 2777 27591 2835 27597
rect 2777 27557 2789 27591
rect 2823 27588 2835 27591
rect 2866 27588 2872 27600
rect 2823 27560 2872 27588
rect 2823 27557 2835 27560
rect 2777 27551 2835 27557
rect 2866 27548 2872 27560
rect 2924 27548 2930 27600
rect 3973 27591 4031 27597
rect 3973 27557 3985 27591
rect 4019 27588 4031 27591
rect 4062 27588 4068 27600
rect 4019 27560 4068 27588
rect 4019 27557 4031 27560
rect 3973 27551 4031 27557
rect 4062 27548 4068 27560
rect 4120 27548 4126 27600
rect 4614 27588 4620 27600
rect 4575 27560 4620 27588
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 5994 27588 6000 27600
rect 5955 27560 6000 27588
rect 5994 27548 6000 27560
rect 6052 27548 6058 27600
rect 7098 27588 7104 27600
rect 7059 27560 7104 27588
rect 7098 27548 7104 27560
rect 7156 27548 7162 27600
rect 8570 27588 8576 27600
rect 8531 27560 8576 27588
rect 8570 27548 8576 27560
rect 8628 27548 8634 27600
rect 9582 27588 9588 27600
rect 9543 27560 9588 27588
rect 9582 27548 9588 27560
rect 9640 27548 9646 27600
rect 11146 27588 11152 27600
rect 11107 27560 11152 27588
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 12066 27588 12072 27600
rect 12027 27560 12072 27588
rect 12066 27548 12072 27560
rect 12124 27548 12130 27600
rect 13814 27548 13820 27600
rect 13872 27588 13878 27600
rect 14277 27591 14335 27597
rect 14277 27588 14289 27591
rect 13872 27560 14289 27588
rect 13872 27548 13878 27560
rect 14277 27557 14289 27560
rect 14323 27557 14335 27591
rect 14918 27588 14924 27600
rect 14879 27560 14924 27588
rect 14277 27551 14335 27557
rect 14918 27548 14924 27560
rect 14976 27548 14982 27600
rect 16574 27548 16580 27600
rect 16632 27588 16638 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 16632 27560 16865 27588
rect 16632 27548 16638 27560
rect 16853 27557 16865 27560
rect 16899 27557 16911 27591
rect 16853 27551 16911 27557
rect 16942 27548 16948 27600
rect 17000 27588 17006 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17000 27560 17509 27588
rect 17000 27548 17006 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 18690 27588 18696 27600
rect 18651 27560 18696 27588
rect 17497 27551 17555 27557
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 19518 27588 19524 27600
rect 19479 27560 19524 27588
rect 19518 27548 19524 27560
rect 19576 27548 19582 27600
rect 21174 27588 21180 27600
rect 21135 27560 21180 27588
rect 21174 27548 21180 27560
rect 21232 27548 21238 27600
rect 22002 27588 22008 27600
rect 21963 27560 22008 27588
rect 22002 27548 22008 27560
rect 22060 27548 22066 27600
rect 1104 27226 22976 27248
rect 1104 27174 6378 27226
rect 6430 27174 6442 27226
rect 6494 27174 6506 27226
rect 6558 27174 6570 27226
rect 6622 27174 6634 27226
rect 6686 27174 11806 27226
rect 11858 27174 11870 27226
rect 11922 27174 11934 27226
rect 11986 27174 11998 27226
rect 12050 27174 12062 27226
rect 12114 27174 17234 27226
rect 17286 27174 17298 27226
rect 17350 27174 17362 27226
rect 17414 27174 17426 27226
rect 17478 27174 17490 27226
rect 17542 27174 22662 27226
rect 22714 27174 22726 27226
rect 22778 27174 22790 27226
rect 22842 27174 22854 27226
rect 22906 27174 22918 27226
rect 22970 27174 22976 27226
rect 1104 27152 22976 27174
rect 1394 26936 1400 26988
rect 1452 26976 1458 26988
rect 1581 26979 1639 26985
rect 1581 26976 1593 26979
rect 1452 26948 1593 26976
rect 1452 26936 1458 26948
rect 1581 26945 1593 26948
rect 1627 26945 1639 26979
rect 1581 26939 1639 26945
rect 2225 26979 2283 26985
rect 2225 26945 2237 26979
rect 2271 26976 2283 26979
rect 2774 26976 2780 26988
rect 2271 26948 2780 26976
rect 2271 26945 2283 26948
rect 2225 26939 2283 26945
rect 2774 26936 2780 26948
rect 2832 26936 2838 26988
rect 22278 26840 22284 26852
rect 22239 26812 22284 26840
rect 22278 26800 22284 26812
rect 22336 26800 22342 26852
rect 1104 26682 22816 26704
rect 1104 26630 3664 26682
rect 3716 26630 3728 26682
rect 3780 26630 3792 26682
rect 3844 26630 3856 26682
rect 3908 26630 3920 26682
rect 3972 26630 9092 26682
rect 9144 26630 9156 26682
rect 9208 26630 9220 26682
rect 9272 26630 9284 26682
rect 9336 26630 9348 26682
rect 9400 26630 14520 26682
rect 14572 26630 14584 26682
rect 14636 26630 14648 26682
rect 14700 26630 14712 26682
rect 14764 26630 14776 26682
rect 14828 26630 19948 26682
rect 20000 26630 20012 26682
rect 20064 26630 20076 26682
rect 20128 26630 20140 26682
rect 20192 26630 20204 26682
rect 20256 26630 22816 26682
rect 1104 26608 22816 26630
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 22278 26364 22284 26376
rect 22239 26336 22284 26364
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 1104 26138 22976 26160
rect 1104 26086 6378 26138
rect 6430 26086 6442 26138
rect 6494 26086 6506 26138
rect 6558 26086 6570 26138
rect 6622 26086 6634 26138
rect 6686 26086 11806 26138
rect 11858 26086 11870 26138
rect 11922 26086 11934 26138
rect 11986 26086 11998 26138
rect 12050 26086 12062 26138
rect 12114 26086 17234 26138
rect 17286 26086 17298 26138
rect 17350 26086 17362 26138
rect 17414 26086 17426 26138
rect 17478 26086 17490 26138
rect 17542 26086 22662 26138
rect 22714 26086 22726 26138
rect 22778 26086 22790 26138
rect 22842 26086 22854 26138
rect 22906 26086 22918 26138
rect 22970 26086 22976 26138
rect 1104 26064 22976 26086
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 1104 25594 22816 25616
rect 1104 25542 3664 25594
rect 3716 25542 3728 25594
rect 3780 25542 3792 25594
rect 3844 25542 3856 25594
rect 3908 25542 3920 25594
rect 3972 25542 9092 25594
rect 9144 25542 9156 25594
rect 9208 25542 9220 25594
rect 9272 25542 9284 25594
rect 9336 25542 9348 25594
rect 9400 25542 14520 25594
rect 14572 25542 14584 25594
rect 14636 25542 14648 25594
rect 14700 25542 14712 25594
rect 14764 25542 14776 25594
rect 14828 25542 19948 25594
rect 20000 25542 20012 25594
rect 20064 25542 20076 25594
rect 20128 25542 20140 25594
rect 20192 25542 20204 25594
rect 20256 25542 22816 25594
rect 1104 25520 22816 25542
rect 22278 25276 22284 25288
rect 22239 25248 22284 25276
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 1104 25050 22976 25072
rect 1104 24998 6378 25050
rect 6430 24998 6442 25050
rect 6494 24998 6506 25050
rect 6558 24998 6570 25050
rect 6622 24998 6634 25050
rect 6686 24998 11806 25050
rect 11858 24998 11870 25050
rect 11922 24998 11934 25050
rect 11986 24998 11998 25050
rect 12050 24998 12062 25050
rect 12114 24998 17234 25050
rect 17286 24998 17298 25050
rect 17350 24998 17362 25050
rect 17414 24998 17426 25050
rect 17478 24998 17490 25050
rect 17542 24998 22662 25050
rect 22714 24998 22726 25050
rect 22778 24998 22790 25050
rect 22842 24998 22854 25050
rect 22906 24998 22918 25050
rect 22970 24998 22976 25050
rect 1104 24976 22976 24998
rect 22278 24664 22284 24676
rect 22239 24636 22284 24664
rect 22278 24624 22284 24636
rect 22336 24624 22342 24676
rect 1104 24506 22816 24528
rect 1104 24454 3664 24506
rect 3716 24454 3728 24506
rect 3780 24454 3792 24506
rect 3844 24454 3856 24506
rect 3908 24454 3920 24506
rect 3972 24454 9092 24506
rect 9144 24454 9156 24506
rect 9208 24454 9220 24506
rect 9272 24454 9284 24506
rect 9336 24454 9348 24506
rect 9400 24454 14520 24506
rect 14572 24454 14584 24506
rect 14636 24454 14648 24506
rect 14700 24454 14712 24506
rect 14764 24454 14776 24506
rect 14828 24454 19948 24506
rect 20000 24454 20012 24506
rect 20064 24454 20076 24506
rect 20128 24454 20140 24506
rect 20192 24454 20204 24506
rect 20256 24454 22816 24506
rect 1104 24432 22816 24454
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 1104 23962 22976 23984
rect 1104 23910 6378 23962
rect 6430 23910 6442 23962
rect 6494 23910 6506 23962
rect 6558 23910 6570 23962
rect 6622 23910 6634 23962
rect 6686 23910 11806 23962
rect 11858 23910 11870 23962
rect 11922 23910 11934 23962
rect 11986 23910 11998 23962
rect 12050 23910 12062 23962
rect 12114 23910 17234 23962
rect 17286 23910 17298 23962
rect 17350 23910 17362 23962
rect 17414 23910 17426 23962
rect 17478 23910 17490 23962
rect 17542 23910 22662 23962
rect 22714 23910 22726 23962
rect 22778 23910 22790 23962
rect 22842 23910 22854 23962
rect 22906 23910 22918 23962
rect 22970 23910 22976 23962
rect 1104 23888 22976 23910
rect 22278 23576 22284 23588
rect 22239 23548 22284 23576
rect 22278 23536 22284 23548
rect 22336 23536 22342 23588
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 1104 23418 22816 23440
rect 1104 23366 3664 23418
rect 3716 23366 3728 23418
rect 3780 23366 3792 23418
rect 3844 23366 3856 23418
rect 3908 23366 3920 23418
rect 3972 23366 9092 23418
rect 9144 23366 9156 23418
rect 9208 23366 9220 23418
rect 9272 23366 9284 23418
rect 9336 23366 9348 23418
rect 9400 23366 14520 23418
rect 14572 23366 14584 23418
rect 14636 23366 14648 23418
rect 14700 23366 14712 23418
rect 14764 23366 14776 23418
rect 14828 23366 19948 23418
rect 20000 23366 20012 23418
rect 20064 23366 20076 23418
rect 20128 23366 20140 23418
rect 20192 23366 20204 23418
rect 20256 23366 22816 23418
rect 1104 23344 22816 23366
rect 22278 23100 22284 23112
rect 22239 23072 22284 23100
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 1104 22874 22976 22896
rect 1104 22822 6378 22874
rect 6430 22822 6442 22874
rect 6494 22822 6506 22874
rect 6558 22822 6570 22874
rect 6622 22822 6634 22874
rect 6686 22822 11806 22874
rect 11858 22822 11870 22874
rect 11922 22822 11934 22874
rect 11986 22822 11998 22874
rect 12050 22822 12062 22874
rect 12114 22822 17234 22874
rect 17286 22822 17298 22874
rect 17350 22822 17362 22874
rect 17414 22822 17426 22874
rect 17478 22822 17490 22874
rect 17542 22822 22662 22874
rect 22714 22822 22726 22874
rect 22778 22822 22790 22874
rect 22842 22822 22854 22874
rect 22906 22822 22918 22874
rect 22970 22822 22976 22874
rect 1104 22800 22976 22822
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 1104 22330 22816 22352
rect 1104 22278 3664 22330
rect 3716 22278 3728 22330
rect 3780 22278 3792 22330
rect 3844 22278 3856 22330
rect 3908 22278 3920 22330
rect 3972 22278 9092 22330
rect 9144 22278 9156 22330
rect 9208 22278 9220 22330
rect 9272 22278 9284 22330
rect 9336 22278 9348 22330
rect 9400 22278 14520 22330
rect 14572 22278 14584 22330
rect 14636 22278 14648 22330
rect 14700 22278 14712 22330
rect 14764 22278 14776 22330
rect 14828 22278 19948 22330
rect 20000 22278 20012 22330
rect 20064 22278 20076 22330
rect 20128 22278 20140 22330
rect 20192 22278 20204 22330
rect 20256 22278 22816 22330
rect 1104 22256 22816 22278
rect 22278 22148 22284 22160
rect 22239 22120 22284 22148
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 1578 21468 1584 21480
rect 1539 21440 1584 21468
rect 1578 21428 1584 21440
rect 1636 21428 1642 21480
rect 22278 21400 22284 21412
rect 22239 21372 22284 21400
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 22278 20312 22284 20324
rect 22239 20284 22284 20312
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 22278 19836 22284 19848
rect 22239 19808 22284 19836
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 22278 18748 22284 18760
rect 22239 18720 22284 18748
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 22278 18136 22284 18148
rect 22239 18108 22284 18136
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 22278 17048 22284 17060
rect 22239 17020 22284 17048
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 22278 16640 22284 16652
rect 22239 16612 22284 16640
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 22278 15484 22284 15496
rect 22239 15456 22284 15484
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 22278 14872 22284 14884
rect 22239 14844 22284 14872
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 22278 13852 22284 13864
rect 22239 13824 22284 13852
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 22278 13308 22284 13320
rect 22239 13280 22284 13308
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 22278 12220 22284 12232
rect 22239 12192 22284 12220
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 22278 11608 22284 11620
rect 22239 11580 22284 11608
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 22278 10520 22284 10532
rect 22239 10492 22284 10520
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 22278 10044 22284 10056
rect 22239 10016 22284 10044
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 22278 8956 22284 8968
rect 22239 8928 22284 8956
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 22278 8344 22284 8356
rect 22239 8316 22284 8344
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 22278 7256 22284 7268
rect 22239 7228 22284 7256
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 22278 6780 22284 6792
rect 22239 6752 22284 6780
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 22278 5692 22284 5704
rect 22239 5664 22284 5692
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 22278 5080 22284 5092
rect 22239 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 22278 3992 22284 4004
rect 22239 3964 22284 3992
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 22278 3516 22284 3528
rect 22239 3488 22284 3516
rect 22278 3476 22284 3488
rect 22336 3476 22342 3528
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 3664 27718 3716 27770
rect 3728 27718 3780 27770
rect 3792 27718 3844 27770
rect 3856 27718 3908 27770
rect 3920 27718 3972 27770
rect 9092 27718 9144 27770
rect 9156 27718 9208 27770
rect 9220 27718 9272 27770
rect 9284 27718 9336 27770
rect 9348 27718 9400 27770
rect 14520 27718 14572 27770
rect 14584 27718 14636 27770
rect 14648 27718 14700 27770
rect 14712 27718 14764 27770
rect 14776 27718 14828 27770
rect 19948 27718 20000 27770
rect 20012 27718 20064 27770
rect 20076 27718 20128 27770
rect 20140 27718 20192 27770
rect 20204 27718 20256 27770
rect 2136 27591 2188 27600
rect 2136 27557 2145 27591
rect 2145 27557 2179 27591
rect 2179 27557 2188 27591
rect 2136 27548 2188 27557
rect 2872 27548 2924 27600
rect 4068 27548 4120 27600
rect 4620 27591 4672 27600
rect 4620 27557 4629 27591
rect 4629 27557 4663 27591
rect 4663 27557 4672 27591
rect 4620 27548 4672 27557
rect 6000 27591 6052 27600
rect 6000 27557 6009 27591
rect 6009 27557 6043 27591
rect 6043 27557 6052 27591
rect 6000 27548 6052 27557
rect 7104 27591 7156 27600
rect 7104 27557 7113 27591
rect 7113 27557 7147 27591
rect 7147 27557 7156 27591
rect 7104 27548 7156 27557
rect 8576 27591 8628 27600
rect 8576 27557 8585 27591
rect 8585 27557 8619 27591
rect 8619 27557 8628 27591
rect 8576 27548 8628 27557
rect 9588 27591 9640 27600
rect 9588 27557 9597 27591
rect 9597 27557 9631 27591
rect 9631 27557 9640 27591
rect 9588 27548 9640 27557
rect 11152 27591 11204 27600
rect 11152 27557 11161 27591
rect 11161 27557 11195 27591
rect 11195 27557 11204 27591
rect 11152 27548 11204 27557
rect 12072 27591 12124 27600
rect 12072 27557 12081 27591
rect 12081 27557 12115 27591
rect 12115 27557 12124 27591
rect 12072 27548 12124 27557
rect 13820 27548 13872 27600
rect 14924 27591 14976 27600
rect 14924 27557 14933 27591
rect 14933 27557 14967 27591
rect 14967 27557 14976 27591
rect 14924 27548 14976 27557
rect 16580 27548 16632 27600
rect 16948 27548 17000 27600
rect 18696 27591 18748 27600
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 19524 27591 19576 27600
rect 19524 27557 19533 27591
rect 19533 27557 19567 27591
rect 19567 27557 19576 27591
rect 19524 27548 19576 27557
rect 21180 27591 21232 27600
rect 21180 27557 21189 27591
rect 21189 27557 21223 27591
rect 21223 27557 21232 27591
rect 21180 27548 21232 27557
rect 22008 27591 22060 27600
rect 22008 27557 22017 27591
rect 22017 27557 22051 27591
rect 22051 27557 22060 27591
rect 22008 27548 22060 27557
rect 6378 27174 6430 27226
rect 6442 27174 6494 27226
rect 6506 27174 6558 27226
rect 6570 27174 6622 27226
rect 6634 27174 6686 27226
rect 11806 27174 11858 27226
rect 11870 27174 11922 27226
rect 11934 27174 11986 27226
rect 11998 27174 12050 27226
rect 12062 27174 12114 27226
rect 17234 27174 17286 27226
rect 17298 27174 17350 27226
rect 17362 27174 17414 27226
rect 17426 27174 17478 27226
rect 17490 27174 17542 27226
rect 22662 27174 22714 27226
rect 22726 27174 22778 27226
rect 22790 27174 22842 27226
rect 22854 27174 22906 27226
rect 22918 27174 22970 27226
rect 1400 26936 1452 26988
rect 2780 26936 2832 26988
rect 22284 26843 22336 26852
rect 22284 26809 22293 26843
rect 22293 26809 22327 26843
rect 22327 26809 22336 26843
rect 22284 26800 22336 26809
rect 3664 26630 3716 26682
rect 3728 26630 3780 26682
rect 3792 26630 3844 26682
rect 3856 26630 3908 26682
rect 3920 26630 3972 26682
rect 9092 26630 9144 26682
rect 9156 26630 9208 26682
rect 9220 26630 9272 26682
rect 9284 26630 9336 26682
rect 9348 26630 9400 26682
rect 14520 26630 14572 26682
rect 14584 26630 14636 26682
rect 14648 26630 14700 26682
rect 14712 26630 14764 26682
rect 14776 26630 14828 26682
rect 19948 26630 20000 26682
rect 20012 26630 20064 26682
rect 20076 26630 20128 26682
rect 20140 26630 20192 26682
rect 20204 26630 20256 26682
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 6378 26086 6430 26138
rect 6442 26086 6494 26138
rect 6506 26086 6558 26138
rect 6570 26086 6622 26138
rect 6634 26086 6686 26138
rect 11806 26086 11858 26138
rect 11870 26086 11922 26138
rect 11934 26086 11986 26138
rect 11998 26086 12050 26138
rect 12062 26086 12114 26138
rect 17234 26086 17286 26138
rect 17298 26086 17350 26138
rect 17362 26086 17414 26138
rect 17426 26086 17478 26138
rect 17490 26086 17542 26138
rect 22662 26086 22714 26138
rect 22726 26086 22778 26138
rect 22790 26086 22842 26138
rect 22854 26086 22906 26138
rect 22918 26086 22970 26138
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 3664 25542 3716 25594
rect 3728 25542 3780 25594
rect 3792 25542 3844 25594
rect 3856 25542 3908 25594
rect 3920 25542 3972 25594
rect 9092 25542 9144 25594
rect 9156 25542 9208 25594
rect 9220 25542 9272 25594
rect 9284 25542 9336 25594
rect 9348 25542 9400 25594
rect 14520 25542 14572 25594
rect 14584 25542 14636 25594
rect 14648 25542 14700 25594
rect 14712 25542 14764 25594
rect 14776 25542 14828 25594
rect 19948 25542 20000 25594
rect 20012 25542 20064 25594
rect 20076 25542 20128 25594
rect 20140 25542 20192 25594
rect 20204 25542 20256 25594
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 22284 25236 22336 25245
rect 6378 24998 6430 25050
rect 6442 24998 6494 25050
rect 6506 24998 6558 25050
rect 6570 24998 6622 25050
rect 6634 24998 6686 25050
rect 11806 24998 11858 25050
rect 11870 24998 11922 25050
rect 11934 24998 11986 25050
rect 11998 24998 12050 25050
rect 12062 24998 12114 25050
rect 17234 24998 17286 25050
rect 17298 24998 17350 25050
rect 17362 24998 17414 25050
rect 17426 24998 17478 25050
rect 17490 24998 17542 25050
rect 22662 24998 22714 25050
rect 22726 24998 22778 25050
rect 22790 24998 22842 25050
rect 22854 24998 22906 25050
rect 22918 24998 22970 25050
rect 22284 24667 22336 24676
rect 22284 24633 22293 24667
rect 22293 24633 22327 24667
rect 22327 24633 22336 24667
rect 22284 24624 22336 24633
rect 3664 24454 3716 24506
rect 3728 24454 3780 24506
rect 3792 24454 3844 24506
rect 3856 24454 3908 24506
rect 3920 24454 3972 24506
rect 9092 24454 9144 24506
rect 9156 24454 9208 24506
rect 9220 24454 9272 24506
rect 9284 24454 9336 24506
rect 9348 24454 9400 24506
rect 14520 24454 14572 24506
rect 14584 24454 14636 24506
rect 14648 24454 14700 24506
rect 14712 24454 14764 24506
rect 14776 24454 14828 24506
rect 19948 24454 20000 24506
rect 20012 24454 20064 24506
rect 20076 24454 20128 24506
rect 20140 24454 20192 24506
rect 20204 24454 20256 24506
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 6378 23910 6430 23962
rect 6442 23910 6494 23962
rect 6506 23910 6558 23962
rect 6570 23910 6622 23962
rect 6634 23910 6686 23962
rect 11806 23910 11858 23962
rect 11870 23910 11922 23962
rect 11934 23910 11986 23962
rect 11998 23910 12050 23962
rect 12062 23910 12114 23962
rect 17234 23910 17286 23962
rect 17298 23910 17350 23962
rect 17362 23910 17414 23962
rect 17426 23910 17478 23962
rect 17490 23910 17542 23962
rect 22662 23910 22714 23962
rect 22726 23910 22778 23962
rect 22790 23910 22842 23962
rect 22854 23910 22906 23962
rect 22918 23910 22970 23962
rect 22284 23579 22336 23588
rect 22284 23545 22293 23579
rect 22293 23545 22327 23579
rect 22327 23545 22336 23579
rect 22284 23536 22336 23545
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 3664 23366 3716 23418
rect 3728 23366 3780 23418
rect 3792 23366 3844 23418
rect 3856 23366 3908 23418
rect 3920 23366 3972 23418
rect 9092 23366 9144 23418
rect 9156 23366 9208 23418
rect 9220 23366 9272 23418
rect 9284 23366 9336 23418
rect 9348 23366 9400 23418
rect 14520 23366 14572 23418
rect 14584 23366 14636 23418
rect 14648 23366 14700 23418
rect 14712 23366 14764 23418
rect 14776 23366 14828 23418
rect 19948 23366 20000 23418
rect 20012 23366 20064 23418
rect 20076 23366 20128 23418
rect 20140 23366 20192 23418
rect 20204 23366 20256 23418
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 6378 22822 6430 22874
rect 6442 22822 6494 22874
rect 6506 22822 6558 22874
rect 6570 22822 6622 22874
rect 6634 22822 6686 22874
rect 11806 22822 11858 22874
rect 11870 22822 11922 22874
rect 11934 22822 11986 22874
rect 11998 22822 12050 22874
rect 12062 22822 12114 22874
rect 17234 22822 17286 22874
rect 17298 22822 17350 22874
rect 17362 22822 17414 22874
rect 17426 22822 17478 22874
rect 17490 22822 17542 22874
rect 22662 22822 22714 22874
rect 22726 22822 22778 22874
rect 22790 22822 22842 22874
rect 22854 22822 22906 22874
rect 22918 22822 22970 22874
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 3664 22278 3716 22330
rect 3728 22278 3780 22330
rect 3792 22278 3844 22330
rect 3856 22278 3908 22330
rect 3920 22278 3972 22330
rect 9092 22278 9144 22330
rect 9156 22278 9208 22330
rect 9220 22278 9272 22330
rect 9284 22278 9336 22330
rect 9348 22278 9400 22330
rect 14520 22278 14572 22330
rect 14584 22278 14636 22330
rect 14648 22278 14700 22330
rect 14712 22278 14764 22330
rect 14776 22278 14828 22330
rect 19948 22278 20000 22330
rect 20012 22278 20064 22330
rect 20076 22278 20128 22330
rect 20140 22278 20192 22330
rect 20204 22278 20256 22330
rect 22284 22151 22336 22160
rect 22284 22117 22293 22151
rect 22293 22117 22327 22151
rect 22327 22117 22336 22151
rect 22284 22108 22336 22117
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 1584 21471 1636 21480
rect 1584 21437 1593 21471
rect 1593 21437 1627 21471
rect 1627 21437 1636 21471
rect 1584 21428 1636 21437
rect 22284 21403 22336 21412
rect 22284 21369 22293 21403
rect 22293 21369 22327 21403
rect 22327 21369 22336 21403
rect 22284 21360 22336 21369
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 22284 20315 22336 20324
rect 22284 20281 22293 20315
rect 22293 20281 22327 20315
rect 22327 20281 22336 20315
rect 22284 20272 22336 20281
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 22284 18139 22336 18148
rect 22284 18105 22293 18139
rect 22293 18105 22327 18139
rect 22327 18105 22336 18139
rect 22284 18096 22336 18105
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 22284 17051 22336 17060
rect 22284 17017 22293 17051
rect 22293 17017 22327 17051
rect 22327 17017 22336 17051
rect 22284 17008 22336 17017
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 22284 14875 22336 14884
rect 22284 14841 22293 14875
rect 22293 14841 22327 14875
rect 22327 14841 22336 14875
rect 22284 14832 22336 14841
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 22284 13311 22336 13320
rect 22284 13277 22293 13311
rect 22293 13277 22327 13311
rect 22327 13277 22336 13311
rect 22284 13268 22336 13277
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 22284 11611 22336 11620
rect 22284 11577 22293 11611
rect 22293 11577 22327 11611
rect 22327 11577 22336 11611
rect 22284 11568 22336 11577
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 22284 10523 22336 10532
rect 22284 10489 22293 10523
rect 22293 10489 22327 10523
rect 22327 10489 22336 10523
rect 22284 10480 22336 10489
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 22284 8347 22336 8356
rect 22284 8313 22293 8347
rect 22293 8313 22327 8347
rect 22327 8313 22336 8347
rect 22284 8304 22336 8313
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 22284 7259 22336 7268
rect 22284 7225 22293 7259
rect 22293 7225 22327 7259
rect 22327 7225 22336 7259
rect 22284 7216 22336 7225
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 22284 6783 22336 6792
rect 22284 6749 22293 6783
rect 22293 6749 22327 6783
rect 22327 6749 22336 6783
rect 22284 6740 22336 6749
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 22284 5083 22336 5092
rect 22284 5049 22293 5083
rect 22293 5049 22327 5083
rect 22327 5049 22336 5083
rect 22284 5040 22336 5049
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 22284 3995 22336 4004
rect 22284 3961 22293 3995
rect 22293 3961 22327 3995
rect 22327 3961 22336 3995
rect 22284 3952 22336 3961
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 22284 3519 22336 3528
rect 22284 3485 22293 3519
rect 22293 3485 22327 3519
rect 22327 3485 22336 3519
rect 22284 3476 22336 3485
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 1400 2796 1452 2848
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 1214 29322 1270 30000
rect 2042 29322 2098 30000
rect 1214 29294 1348 29322
rect 1214 29200 1270 29294
rect 1320 27010 1348 29294
rect 2042 29294 2176 29322
rect 2042 29200 2098 29294
rect 2148 27606 2176 29294
rect 2870 29200 2926 30000
rect 3698 29322 3754 30000
rect 4526 29322 4582 30000
rect 3698 29294 4108 29322
rect 3698 29200 3754 29294
rect 2870 28248 2926 28257
rect 2870 28183 2926 28192
rect 2884 27606 2912 28183
rect 3664 27772 3972 27781
rect 3664 27770 3670 27772
rect 3726 27770 3750 27772
rect 3806 27770 3830 27772
rect 3886 27770 3910 27772
rect 3966 27770 3972 27772
rect 3726 27718 3728 27770
rect 3908 27718 3910 27770
rect 3664 27716 3670 27718
rect 3726 27716 3750 27718
rect 3806 27716 3830 27718
rect 3886 27716 3910 27718
rect 3966 27716 3972 27718
rect 3664 27707 3972 27716
rect 4080 27606 4108 29294
rect 4526 29294 4660 29322
rect 4526 29200 4582 29294
rect 4632 27606 4660 29294
rect 5354 29200 5410 30000
rect 6182 29322 6238 30000
rect 6012 29294 6238 29322
rect 6012 27606 6040 29294
rect 6182 29200 6238 29294
rect 7010 29322 7066 30000
rect 7010 29294 7144 29322
rect 7010 29200 7066 29294
rect 7116 27606 7144 29294
rect 7838 29200 7894 30000
rect 8666 29322 8722 30000
rect 8588 29294 8722 29322
rect 8588 27606 8616 29294
rect 8666 29200 8722 29294
rect 9494 29322 9550 30000
rect 9494 29294 9628 29322
rect 9494 29200 9550 29294
rect 9092 27772 9400 27781
rect 9092 27770 9098 27772
rect 9154 27770 9178 27772
rect 9234 27770 9258 27772
rect 9314 27770 9338 27772
rect 9394 27770 9400 27772
rect 9154 27718 9156 27770
rect 9336 27718 9338 27770
rect 9092 27716 9098 27718
rect 9154 27716 9178 27718
rect 9234 27716 9258 27718
rect 9314 27716 9338 27718
rect 9394 27716 9400 27718
rect 9092 27707 9400 27716
rect 9600 27606 9628 29294
rect 10322 29200 10378 30000
rect 11150 29200 11206 30000
rect 11978 29322 12034 30000
rect 11978 29294 12112 29322
rect 11978 29200 12034 29294
rect 11164 27606 11192 29200
rect 12084 27606 12112 29294
rect 12806 29200 12862 30000
rect 13634 29322 13690 30000
rect 14462 29322 14518 30000
rect 13634 29294 13768 29322
rect 13634 29200 13690 29294
rect 2136 27600 2188 27606
rect 2872 27600 2924 27606
rect 2136 27542 2188 27548
rect 2778 27568 2834 27577
rect 2872 27542 2924 27548
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 6000 27600 6052 27606
rect 6000 27542 6052 27548
rect 7104 27600 7156 27606
rect 7104 27542 7156 27548
rect 8576 27600 8628 27606
rect 8576 27542 8628 27548
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 12072 27600 12124 27606
rect 13740 27588 13768 29294
rect 14462 29294 14964 29322
rect 14462 29200 14518 29294
rect 14520 27772 14828 27781
rect 14520 27770 14526 27772
rect 14582 27770 14606 27772
rect 14662 27770 14686 27772
rect 14742 27770 14766 27772
rect 14822 27770 14828 27772
rect 14582 27718 14584 27770
rect 14764 27718 14766 27770
rect 14520 27716 14526 27718
rect 14582 27716 14606 27718
rect 14662 27716 14686 27718
rect 14742 27716 14766 27718
rect 14822 27716 14828 27718
rect 14520 27707 14828 27716
rect 14936 27606 14964 29294
rect 15290 29200 15346 30000
rect 16118 29322 16174 30000
rect 16118 29294 16528 29322
rect 16118 29200 16174 29294
rect 13820 27600 13872 27606
rect 13740 27560 13820 27588
rect 12072 27542 12124 27548
rect 13820 27542 13872 27548
rect 14924 27600 14976 27606
rect 16500 27588 16528 29294
rect 16946 29200 17002 30000
rect 17774 29200 17830 30000
rect 18602 29322 18658 30000
rect 19430 29322 19486 30000
rect 18602 29294 18736 29322
rect 18602 29200 18658 29294
rect 16960 27606 16988 29200
rect 18708 27606 18736 29294
rect 19430 29294 19564 29322
rect 19430 29200 19486 29294
rect 19536 27606 19564 29294
rect 20258 29200 20314 30000
rect 21086 29322 21142 30000
rect 21914 29322 21970 30000
rect 21086 29294 21220 29322
rect 21086 29200 21142 29294
rect 19948 27772 20256 27781
rect 19948 27770 19954 27772
rect 20010 27770 20034 27772
rect 20090 27770 20114 27772
rect 20170 27770 20194 27772
rect 20250 27770 20256 27772
rect 20010 27718 20012 27770
rect 20192 27718 20194 27770
rect 19948 27716 19954 27718
rect 20010 27716 20034 27718
rect 20090 27716 20114 27718
rect 20170 27716 20194 27718
rect 20250 27716 20256 27718
rect 19948 27707 20256 27716
rect 21192 27606 21220 29294
rect 21914 29294 22048 29322
rect 21914 29200 21970 29294
rect 22020 27606 22048 29294
rect 22742 29200 22798 30000
rect 16580 27600 16632 27606
rect 16500 27560 16580 27588
rect 14924 27542 14976 27548
rect 16580 27542 16632 27548
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 21180 27600 21232 27606
rect 21180 27542 21232 27548
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 2778 27503 2834 27512
rect 1320 26994 1440 27010
rect 2792 26994 2820 27503
rect 6378 27228 6686 27237
rect 6378 27226 6384 27228
rect 6440 27226 6464 27228
rect 6520 27226 6544 27228
rect 6600 27226 6624 27228
rect 6680 27226 6686 27228
rect 6440 27174 6442 27226
rect 6622 27174 6624 27226
rect 6378 27172 6384 27174
rect 6440 27172 6464 27174
rect 6520 27172 6544 27174
rect 6600 27172 6624 27174
rect 6680 27172 6686 27174
rect 6378 27163 6686 27172
rect 11806 27228 12114 27237
rect 11806 27226 11812 27228
rect 11868 27226 11892 27228
rect 11948 27226 11972 27228
rect 12028 27226 12052 27228
rect 12108 27226 12114 27228
rect 11868 27174 11870 27226
rect 12050 27174 12052 27226
rect 11806 27172 11812 27174
rect 11868 27172 11892 27174
rect 11948 27172 11972 27174
rect 12028 27172 12052 27174
rect 12108 27172 12114 27174
rect 11806 27163 12114 27172
rect 17234 27228 17542 27237
rect 17234 27226 17240 27228
rect 17296 27226 17320 27228
rect 17376 27226 17400 27228
rect 17456 27226 17480 27228
rect 17536 27226 17542 27228
rect 17296 27174 17298 27226
rect 17478 27174 17480 27226
rect 17234 27172 17240 27174
rect 17296 27172 17320 27174
rect 17376 27172 17400 27174
rect 17456 27172 17480 27174
rect 17536 27172 17542 27174
rect 17234 27163 17542 27172
rect 22662 27228 22970 27237
rect 22662 27226 22668 27228
rect 22724 27226 22748 27228
rect 22804 27226 22828 27228
rect 22884 27226 22908 27228
rect 22964 27226 22970 27228
rect 22724 27174 22726 27226
rect 22906 27174 22908 27226
rect 22662 27172 22668 27174
rect 22724 27172 22748 27174
rect 22804 27172 22828 27174
rect 22884 27172 22908 27174
rect 22964 27172 22970 27174
rect 22662 27163 22970 27172
rect 1320 26988 1452 26994
rect 1320 26982 1400 26988
rect 1400 26930 1452 26936
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 22282 26888 22338 26897
rect 22282 26823 22284 26832
rect 22336 26823 22338 26832
rect 22284 26794 22336 26800
rect 3664 26684 3972 26693
rect 3664 26682 3670 26684
rect 3726 26682 3750 26684
rect 3806 26682 3830 26684
rect 3886 26682 3910 26684
rect 3966 26682 3972 26684
rect 3726 26630 3728 26682
rect 3908 26630 3910 26682
rect 3664 26628 3670 26630
rect 3726 26628 3750 26630
rect 3806 26628 3830 26630
rect 3886 26628 3910 26630
rect 3966 26628 3972 26630
rect 3664 26619 3972 26628
rect 9092 26684 9400 26693
rect 9092 26682 9098 26684
rect 9154 26682 9178 26684
rect 9234 26682 9258 26684
rect 9314 26682 9338 26684
rect 9394 26682 9400 26684
rect 9154 26630 9156 26682
rect 9336 26630 9338 26682
rect 9092 26628 9098 26630
rect 9154 26628 9178 26630
rect 9234 26628 9258 26630
rect 9314 26628 9338 26630
rect 9394 26628 9400 26630
rect 9092 26619 9400 26628
rect 14520 26684 14828 26693
rect 14520 26682 14526 26684
rect 14582 26682 14606 26684
rect 14662 26682 14686 26684
rect 14742 26682 14766 26684
rect 14822 26682 14828 26684
rect 14582 26630 14584 26682
rect 14764 26630 14766 26682
rect 14520 26628 14526 26630
rect 14582 26628 14606 26630
rect 14662 26628 14686 26630
rect 14742 26628 14766 26630
rect 14822 26628 14828 26630
rect 14520 26619 14828 26628
rect 19948 26684 20256 26693
rect 19948 26682 19954 26684
rect 20010 26682 20034 26684
rect 20090 26682 20114 26684
rect 20170 26682 20194 26684
rect 20250 26682 20256 26684
rect 20010 26630 20012 26682
rect 20192 26630 20194 26682
rect 19948 26628 19954 26630
rect 20010 26628 20034 26630
rect 20090 26628 20114 26630
rect 20170 26628 20194 26630
rect 20250 26628 20256 26630
rect 19948 26619 20256 26628
rect 1584 26376 1636 26382
rect 22284 26376 22336 26382
rect 1584 26318 1636 26324
rect 22282 26344 22284 26353
rect 22336 26344 22338 26353
rect 1596 26217 1624 26318
rect 22282 26279 22338 26288
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 6378 26140 6686 26149
rect 6378 26138 6384 26140
rect 6440 26138 6464 26140
rect 6520 26138 6544 26140
rect 6600 26138 6624 26140
rect 6680 26138 6686 26140
rect 6440 26086 6442 26138
rect 6622 26086 6624 26138
rect 6378 26084 6384 26086
rect 6440 26084 6464 26086
rect 6520 26084 6544 26086
rect 6600 26084 6624 26086
rect 6680 26084 6686 26086
rect 6378 26075 6686 26084
rect 11806 26140 12114 26149
rect 11806 26138 11812 26140
rect 11868 26138 11892 26140
rect 11948 26138 11972 26140
rect 12028 26138 12052 26140
rect 12108 26138 12114 26140
rect 11868 26086 11870 26138
rect 12050 26086 12052 26138
rect 11806 26084 11812 26086
rect 11868 26084 11892 26086
rect 11948 26084 11972 26086
rect 12028 26084 12052 26086
rect 12108 26084 12114 26086
rect 11806 26075 12114 26084
rect 17234 26140 17542 26149
rect 17234 26138 17240 26140
rect 17296 26138 17320 26140
rect 17376 26138 17400 26140
rect 17456 26138 17480 26140
rect 17536 26138 17542 26140
rect 17296 26086 17298 26138
rect 17478 26086 17480 26138
rect 17234 26084 17240 26086
rect 17296 26084 17320 26086
rect 17376 26084 17400 26086
rect 17456 26084 17480 26086
rect 17536 26084 17542 26086
rect 17234 26075 17542 26084
rect 22662 26140 22970 26149
rect 22662 26138 22668 26140
rect 22724 26138 22748 26140
rect 22804 26138 22828 26140
rect 22884 26138 22908 26140
rect 22964 26138 22970 26140
rect 22724 26086 22726 26138
rect 22906 26086 22908 26138
rect 22662 26084 22668 26086
rect 22724 26084 22748 26086
rect 22804 26084 22828 26086
rect 22884 26084 22908 26086
rect 22964 26084 22970 26086
rect 22662 26075 22970 26084
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25537 1624 25638
rect 3664 25596 3972 25605
rect 3664 25594 3670 25596
rect 3726 25594 3750 25596
rect 3806 25594 3830 25596
rect 3886 25594 3910 25596
rect 3966 25594 3972 25596
rect 3726 25542 3728 25594
rect 3908 25542 3910 25594
rect 3664 25540 3670 25542
rect 3726 25540 3750 25542
rect 3806 25540 3830 25542
rect 3886 25540 3910 25542
rect 3966 25540 3972 25542
rect 1582 25528 1638 25537
rect 3664 25531 3972 25540
rect 9092 25596 9400 25605
rect 9092 25594 9098 25596
rect 9154 25594 9178 25596
rect 9234 25594 9258 25596
rect 9314 25594 9338 25596
rect 9394 25594 9400 25596
rect 9154 25542 9156 25594
rect 9336 25542 9338 25594
rect 9092 25540 9098 25542
rect 9154 25540 9178 25542
rect 9234 25540 9258 25542
rect 9314 25540 9338 25542
rect 9394 25540 9400 25542
rect 9092 25531 9400 25540
rect 14520 25596 14828 25605
rect 14520 25594 14526 25596
rect 14582 25594 14606 25596
rect 14662 25594 14686 25596
rect 14742 25594 14766 25596
rect 14822 25594 14828 25596
rect 14582 25542 14584 25594
rect 14764 25542 14766 25594
rect 14520 25540 14526 25542
rect 14582 25540 14606 25542
rect 14662 25540 14686 25542
rect 14742 25540 14766 25542
rect 14822 25540 14828 25542
rect 14520 25531 14828 25540
rect 19948 25596 20256 25605
rect 19948 25594 19954 25596
rect 20010 25594 20034 25596
rect 20090 25594 20114 25596
rect 20170 25594 20194 25596
rect 20250 25594 20256 25596
rect 20010 25542 20012 25594
rect 20192 25542 20194 25594
rect 19948 25540 19954 25542
rect 20010 25540 20034 25542
rect 20090 25540 20114 25542
rect 20170 25540 20194 25542
rect 20250 25540 20256 25542
rect 19948 25531 20256 25540
rect 1582 25463 1638 25472
rect 22284 25288 22336 25294
rect 22282 25256 22284 25265
rect 22336 25256 22338 25265
rect 22282 25191 22338 25200
rect 6378 25052 6686 25061
rect 6378 25050 6384 25052
rect 6440 25050 6464 25052
rect 6520 25050 6544 25052
rect 6600 25050 6624 25052
rect 6680 25050 6686 25052
rect 6440 24998 6442 25050
rect 6622 24998 6624 25050
rect 6378 24996 6384 24998
rect 6440 24996 6464 24998
rect 6520 24996 6544 24998
rect 6600 24996 6624 24998
rect 6680 24996 6686 24998
rect 6378 24987 6686 24996
rect 11806 25052 12114 25061
rect 11806 25050 11812 25052
rect 11868 25050 11892 25052
rect 11948 25050 11972 25052
rect 12028 25050 12052 25052
rect 12108 25050 12114 25052
rect 11868 24998 11870 25050
rect 12050 24998 12052 25050
rect 11806 24996 11812 24998
rect 11868 24996 11892 24998
rect 11948 24996 11972 24998
rect 12028 24996 12052 24998
rect 12108 24996 12114 24998
rect 11806 24987 12114 24996
rect 17234 25052 17542 25061
rect 17234 25050 17240 25052
rect 17296 25050 17320 25052
rect 17376 25050 17400 25052
rect 17456 25050 17480 25052
rect 17536 25050 17542 25052
rect 17296 24998 17298 25050
rect 17478 24998 17480 25050
rect 17234 24996 17240 24998
rect 17296 24996 17320 24998
rect 17376 24996 17400 24998
rect 17456 24996 17480 24998
rect 17536 24996 17542 24998
rect 17234 24987 17542 24996
rect 22662 25052 22970 25061
rect 22662 25050 22668 25052
rect 22724 25050 22748 25052
rect 22804 25050 22828 25052
rect 22884 25050 22908 25052
rect 22964 25050 22970 25052
rect 22724 24998 22726 25050
rect 22906 24998 22908 25050
rect 22662 24996 22668 24998
rect 22724 24996 22748 24998
rect 22804 24996 22828 24998
rect 22884 24996 22908 24998
rect 22964 24996 22970 24998
rect 22662 24987 22970 24996
rect 22282 24712 22338 24721
rect 22282 24647 22284 24656
rect 22336 24647 22338 24656
rect 22284 24618 22336 24624
rect 3664 24508 3972 24517
rect 3664 24506 3670 24508
rect 3726 24506 3750 24508
rect 3806 24506 3830 24508
rect 3886 24506 3910 24508
rect 3966 24506 3972 24508
rect 3726 24454 3728 24506
rect 3908 24454 3910 24506
rect 3664 24452 3670 24454
rect 3726 24452 3750 24454
rect 3806 24452 3830 24454
rect 3886 24452 3910 24454
rect 3966 24452 3972 24454
rect 3664 24443 3972 24452
rect 9092 24508 9400 24517
rect 9092 24506 9098 24508
rect 9154 24506 9178 24508
rect 9234 24506 9258 24508
rect 9314 24506 9338 24508
rect 9394 24506 9400 24508
rect 9154 24454 9156 24506
rect 9336 24454 9338 24506
rect 9092 24452 9098 24454
rect 9154 24452 9178 24454
rect 9234 24452 9258 24454
rect 9314 24452 9338 24454
rect 9394 24452 9400 24454
rect 9092 24443 9400 24452
rect 14520 24508 14828 24517
rect 14520 24506 14526 24508
rect 14582 24506 14606 24508
rect 14662 24506 14686 24508
rect 14742 24506 14766 24508
rect 14822 24506 14828 24508
rect 14582 24454 14584 24506
rect 14764 24454 14766 24506
rect 14520 24452 14526 24454
rect 14582 24452 14606 24454
rect 14662 24452 14686 24454
rect 14742 24452 14766 24454
rect 14822 24452 14828 24454
rect 14520 24443 14828 24452
rect 19948 24508 20256 24517
rect 19948 24506 19954 24508
rect 20010 24506 20034 24508
rect 20090 24506 20114 24508
rect 20170 24506 20194 24508
rect 20250 24506 20256 24508
rect 20010 24454 20012 24506
rect 20192 24454 20194 24506
rect 19948 24452 19954 24454
rect 20010 24452 20034 24454
rect 20090 24452 20114 24454
rect 20170 24452 20194 24454
rect 20250 24452 20256 24454
rect 19948 24443 20256 24452
rect 1584 24200 1636 24206
rect 1582 24168 1584 24177
rect 1636 24168 1638 24177
rect 1582 24103 1638 24112
rect 6378 23964 6686 23973
rect 6378 23962 6384 23964
rect 6440 23962 6464 23964
rect 6520 23962 6544 23964
rect 6600 23962 6624 23964
rect 6680 23962 6686 23964
rect 6440 23910 6442 23962
rect 6622 23910 6624 23962
rect 6378 23908 6384 23910
rect 6440 23908 6464 23910
rect 6520 23908 6544 23910
rect 6600 23908 6624 23910
rect 6680 23908 6686 23910
rect 6378 23899 6686 23908
rect 11806 23964 12114 23973
rect 11806 23962 11812 23964
rect 11868 23962 11892 23964
rect 11948 23962 11972 23964
rect 12028 23962 12052 23964
rect 12108 23962 12114 23964
rect 11868 23910 11870 23962
rect 12050 23910 12052 23962
rect 11806 23908 11812 23910
rect 11868 23908 11892 23910
rect 11948 23908 11972 23910
rect 12028 23908 12052 23910
rect 12108 23908 12114 23910
rect 11806 23899 12114 23908
rect 17234 23964 17542 23973
rect 17234 23962 17240 23964
rect 17296 23962 17320 23964
rect 17376 23962 17400 23964
rect 17456 23962 17480 23964
rect 17536 23962 17542 23964
rect 17296 23910 17298 23962
rect 17478 23910 17480 23962
rect 17234 23908 17240 23910
rect 17296 23908 17320 23910
rect 17376 23908 17400 23910
rect 17456 23908 17480 23910
rect 17536 23908 17542 23910
rect 17234 23899 17542 23908
rect 22662 23964 22970 23973
rect 22662 23962 22668 23964
rect 22724 23962 22748 23964
rect 22804 23962 22828 23964
rect 22884 23962 22908 23964
rect 22964 23962 22970 23964
rect 22724 23910 22726 23962
rect 22906 23910 22908 23962
rect 22662 23908 22668 23910
rect 22724 23908 22748 23910
rect 22804 23908 22828 23910
rect 22884 23908 22908 23910
rect 22964 23908 22970 23910
rect 22662 23899 22970 23908
rect 22282 23624 22338 23633
rect 22282 23559 22284 23568
rect 22336 23559 22338 23568
rect 22284 23530 22336 23536
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 3664 23420 3972 23429
rect 3664 23418 3670 23420
rect 3726 23418 3750 23420
rect 3806 23418 3830 23420
rect 3886 23418 3910 23420
rect 3966 23418 3972 23420
rect 3726 23366 3728 23418
rect 3908 23366 3910 23418
rect 3664 23364 3670 23366
rect 3726 23364 3750 23366
rect 3806 23364 3830 23366
rect 3886 23364 3910 23366
rect 3966 23364 3972 23366
rect 3664 23355 3972 23364
rect 9092 23420 9400 23429
rect 9092 23418 9098 23420
rect 9154 23418 9178 23420
rect 9234 23418 9258 23420
rect 9314 23418 9338 23420
rect 9394 23418 9400 23420
rect 9154 23366 9156 23418
rect 9336 23366 9338 23418
rect 9092 23364 9098 23366
rect 9154 23364 9178 23366
rect 9234 23364 9258 23366
rect 9314 23364 9338 23366
rect 9394 23364 9400 23366
rect 9092 23355 9400 23364
rect 14520 23420 14828 23429
rect 14520 23418 14526 23420
rect 14582 23418 14606 23420
rect 14662 23418 14686 23420
rect 14742 23418 14766 23420
rect 14822 23418 14828 23420
rect 14582 23366 14584 23418
rect 14764 23366 14766 23418
rect 14520 23364 14526 23366
rect 14582 23364 14606 23366
rect 14662 23364 14686 23366
rect 14742 23364 14766 23366
rect 14822 23364 14828 23366
rect 14520 23355 14828 23364
rect 19948 23420 20256 23429
rect 19948 23418 19954 23420
rect 20010 23418 20034 23420
rect 20090 23418 20114 23420
rect 20170 23418 20194 23420
rect 20250 23418 20256 23420
rect 20010 23366 20012 23418
rect 20192 23366 20194 23418
rect 19948 23364 19954 23366
rect 20010 23364 20034 23366
rect 20090 23364 20114 23366
rect 20170 23364 20194 23366
rect 20250 23364 20256 23366
rect 19948 23355 20256 23364
rect 22284 23112 22336 23118
rect 22282 23080 22284 23089
rect 22336 23080 22338 23089
rect 22282 23015 22338 23024
rect 6378 22876 6686 22885
rect 6378 22874 6384 22876
rect 6440 22874 6464 22876
rect 6520 22874 6544 22876
rect 6600 22874 6624 22876
rect 6680 22874 6686 22876
rect 6440 22822 6442 22874
rect 6622 22822 6624 22874
rect 6378 22820 6384 22822
rect 6440 22820 6464 22822
rect 6520 22820 6544 22822
rect 6600 22820 6624 22822
rect 6680 22820 6686 22822
rect 6378 22811 6686 22820
rect 11806 22876 12114 22885
rect 11806 22874 11812 22876
rect 11868 22874 11892 22876
rect 11948 22874 11972 22876
rect 12028 22874 12052 22876
rect 12108 22874 12114 22876
rect 11868 22822 11870 22874
rect 12050 22822 12052 22874
rect 11806 22820 11812 22822
rect 11868 22820 11892 22822
rect 11948 22820 11972 22822
rect 12028 22820 12052 22822
rect 12108 22820 12114 22822
rect 11806 22811 12114 22820
rect 17234 22876 17542 22885
rect 17234 22874 17240 22876
rect 17296 22874 17320 22876
rect 17376 22874 17400 22876
rect 17456 22874 17480 22876
rect 17536 22874 17542 22876
rect 17296 22822 17298 22874
rect 17478 22822 17480 22874
rect 17234 22820 17240 22822
rect 17296 22820 17320 22822
rect 17376 22820 17400 22822
rect 17456 22820 17480 22822
rect 17536 22820 17542 22822
rect 17234 22811 17542 22820
rect 22662 22876 22970 22885
rect 22662 22874 22668 22876
rect 22724 22874 22748 22876
rect 22804 22874 22828 22876
rect 22884 22874 22908 22876
rect 22964 22874 22970 22876
rect 22724 22822 22726 22874
rect 22906 22822 22908 22874
rect 22662 22820 22668 22822
rect 22724 22820 22748 22822
rect 22804 22820 22828 22822
rect 22884 22820 22908 22822
rect 22964 22820 22970 22822
rect 22662 22811 22970 22820
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 3664 22332 3972 22341
rect 3664 22330 3670 22332
rect 3726 22330 3750 22332
rect 3806 22330 3830 22332
rect 3886 22330 3910 22332
rect 3966 22330 3972 22332
rect 3726 22278 3728 22330
rect 3908 22278 3910 22330
rect 3664 22276 3670 22278
rect 3726 22276 3750 22278
rect 3806 22276 3830 22278
rect 3886 22276 3910 22278
rect 3966 22276 3972 22278
rect 3664 22267 3972 22276
rect 9092 22332 9400 22341
rect 9092 22330 9098 22332
rect 9154 22330 9178 22332
rect 9234 22330 9258 22332
rect 9314 22330 9338 22332
rect 9394 22330 9400 22332
rect 9154 22278 9156 22330
rect 9336 22278 9338 22330
rect 9092 22276 9098 22278
rect 9154 22276 9178 22278
rect 9234 22276 9258 22278
rect 9314 22276 9338 22278
rect 9394 22276 9400 22278
rect 9092 22267 9400 22276
rect 14520 22332 14828 22341
rect 14520 22330 14526 22332
rect 14582 22330 14606 22332
rect 14662 22330 14686 22332
rect 14742 22330 14766 22332
rect 14822 22330 14828 22332
rect 14582 22278 14584 22330
rect 14764 22278 14766 22330
rect 14520 22276 14526 22278
rect 14582 22276 14606 22278
rect 14662 22276 14686 22278
rect 14742 22276 14766 22278
rect 14822 22276 14828 22278
rect 14520 22267 14828 22276
rect 19948 22332 20256 22341
rect 19948 22330 19954 22332
rect 20010 22330 20034 22332
rect 20090 22330 20114 22332
rect 20170 22330 20194 22332
rect 20250 22330 20256 22332
rect 20010 22278 20012 22330
rect 20192 22278 20194 22330
rect 19948 22276 19954 22278
rect 20010 22276 20034 22278
rect 20090 22276 20114 22278
rect 20170 22276 20194 22278
rect 20250 22276 20256 22278
rect 19948 22267 20256 22276
rect 22284 22160 22336 22166
rect 1582 22128 1638 22137
rect 22284 22102 22336 22108
rect 1582 22063 1638 22072
rect 22296 22001 22324 22102
rect 22282 21992 22338 22001
rect 22282 21927 22338 21936
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 1584 21480 1636 21486
rect 1582 21448 1584 21457
rect 1636 21448 1638 21457
rect 1582 21383 1638 21392
rect 22282 21448 22338 21457
rect 22282 21383 22284 21392
rect 22336 21383 22338 21392
rect 22284 21354 22336 21360
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 22282 20360 22338 20369
rect 22282 20295 22284 20304
rect 22336 20295 22338 20304
rect 22284 20266 22336 20272
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 1582 20088 1638 20097
rect 3664 20091 3972 20100
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 1582 20023 1638 20032
rect 1584 19848 1636 19854
rect 22284 19848 22336 19854
rect 1584 19790 1636 19796
rect 22282 19816 22284 19825
rect 22336 19816 22338 19825
rect 1596 19417 1624 19790
rect 22282 19751 22338 19760
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 22284 18760 22336 18766
rect 22282 18728 22284 18737
rect 22336 18728 22338 18737
rect 22282 18663 22338 18672
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 22282 18184 22338 18193
rect 22282 18119 22284 18128
rect 22336 18119 22338 18128
rect 22284 18090 22336 18096
rect 1584 18080 1636 18086
rect 1582 18048 1584 18057
rect 1636 18048 1638 18057
rect 1582 17983 1638 17992
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17377 1624 17614
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 1582 17368 1638 17377
rect 6378 17371 6686 17380
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 1582 17303 1638 17312
rect 22282 17096 22338 17105
rect 22282 17031 22284 17040
rect 22336 17031 22338 17040
rect 22284 17002 22336 17008
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22296 16561 22324 16594
rect 22282 16552 22338 16561
rect 22282 16487 22338 16496
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 1584 16040 1636 16046
rect 1582 16008 1584 16017
rect 1636 16008 1638 16017
rect 1582 15943 1638 15952
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 1584 15496 1636 15502
rect 22284 15496 22336 15502
rect 1584 15438 1636 15444
rect 22282 15464 22284 15473
rect 22336 15464 22338 15473
rect 1596 15337 1624 15438
rect 22282 15399 22338 15408
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 22282 14920 22338 14929
rect 22282 14855 22284 14864
rect 22336 14855 22338 14864
rect 22284 14826 22336 14832
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 22284 13864 22336 13870
rect 22282 13832 22284 13841
rect 22336 13832 22338 13841
rect 22282 13767 22338 13776
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 1584 13320 1636 13326
rect 1582 13288 1584 13297
rect 22284 13320 22336 13326
rect 1636 13288 1638 13297
rect 1582 13223 1638 13232
rect 22282 13288 22284 13297
rect 22336 13288 22338 13297
rect 22282 13223 22338 13232
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 1584 12232 1636 12238
rect 22284 12232 22336 12238
rect 1584 12174 1636 12180
rect 22282 12200 22284 12209
rect 22336 12200 22338 12209
rect 1596 11937 1624 12174
rect 22282 12135 22338 12144
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 1582 11928 1638 11937
rect 6378 11931 6686 11940
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 1582 11863 1638 11872
rect 22282 11656 22338 11665
rect 22282 11591 22284 11600
rect 22336 11591 22338 11600
rect 22284 11562 22336 11568
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11257 1624 11494
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 22282 10568 22338 10577
rect 22282 10503 22284 10512
rect 22336 10503 22338 10512
rect 22284 10474 22336 10480
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 1584 10056 1636 10062
rect 22284 10056 22336 10062
rect 1584 9998 1636 10004
rect 22282 10024 22284 10033
rect 22336 10024 22338 10033
rect 1596 9897 1624 9998
rect 22282 9959 22338 9968
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 1582 9208 1638 9217
rect 3664 9211 3972 9220
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 1582 9143 1638 9152
rect 22284 8968 22336 8974
rect 22282 8936 22284 8945
rect 22336 8936 22338 8945
rect 22282 8871 22338 8880
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 22282 8392 22338 8401
rect 22282 8327 22284 8336
rect 22336 8327 22338 8336
rect 22284 8298 22336 8304
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 1584 7880 1636 7886
rect 1582 7848 1584 7857
rect 1636 7848 1638 7857
rect 1582 7783 1638 7792
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 22282 7304 22338 7313
rect 22282 7239 22284 7248
rect 22336 7239 22338 7248
rect 22284 7210 22336 7216
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 22284 6792 22336 6798
rect 22282 6760 22284 6769
rect 22336 6760 22338 6769
rect 22282 6695 22338 6704
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5817 1624 6054
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 22284 5704 22336 5710
rect 22282 5672 22284 5681
rect 22336 5672 22338 5681
rect 22282 5607 22338 5616
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 1584 5160 1636 5166
rect 1582 5128 1584 5137
rect 1636 5128 1638 5137
rect 1582 5063 1638 5072
rect 22282 5128 22338 5137
rect 22282 5063 22284 5072
rect 22336 5063 22338 5072
rect 22284 5034 22336 5040
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 22282 4040 22338 4049
rect 22282 3975 22284 3984
rect 22336 3975 22338 3984
rect 22284 3946 22336 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3777 1624 3878
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 1582 3768 1638 3777
rect 3664 3771 3972 3780
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 1582 3703 1638 3712
rect 1584 3528 1636 3534
rect 22284 3528 22336 3534
rect 1584 3470 1636 3476
rect 22282 3496 22284 3505
rect 22336 3496 22338 3505
rect 1596 3097 1624 3470
rect 22282 3431 22338 3440
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 1057 1440 2790
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1596 1737 1624 2382
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
rect 1582 1728 1638 1737
rect 1582 1663 1638 1672
rect 1398 1048 1454 1057
rect 1398 983 1454 992
<< via2 >>
rect 2870 28192 2926 28248
rect 3670 27770 3726 27772
rect 3750 27770 3806 27772
rect 3830 27770 3886 27772
rect 3910 27770 3966 27772
rect 3670 27718 3716 27770
rect 3716 27718 3726 27770
rect 3750 27718 3780 27770
rect 3780 27718 3792 27770
rect 3792 27718 3806 27770
rect 3830 27718 3844 27770
rect 3844 27718 3856 27770
rect 3856 27718 3886 27770
rect 3910 27718 3920 27770
rect 3920 27718 3966 27770
rect 3670 27716 3726 27718
rect 3750 27716 3806 27718
rect 3830 27716 3886 27718
rect 3910 27716 3966 27718
rect 9098 27770 9154 27772
rect 9178 27770 9234 27772
rect 9258 27770 9314 27772
rect 9338 27770 9394 27772
rect 9098 27718 9144 27770
rect 9144 27718 9154 27770
rect 9178 27718 9208 27770
rect 9208 27718 9220 27770
rect 9220 27718 9234 27770
rect 9258 27718 9272 27770
rect 9272 27718 9284 27770
rect 9284 27718 9314 27770
rect 9338 27718 9348 27770
rect 9348 27718 9394 27770
rect 9098 27716 9154 27718
rect 9178 27716 9234 27718
rect 9258 27716 9314 27718
rect 9338 27716 9394 27718
rect 2778 27512 2834 27568
rect 14526 27770 14582 27772
rect 14606 27770 14662 27772
rect 14686 27770 14742 27772
rect 14766 27770 14822 27772
rect 14526 27718 14572 27770
rect 14572 27718 14582 27770
rect 14606 27718 14636 27770
rect 14636 27718 14648 27770
rect 14648 27718 14662 27770
rect 14686 27718 14700 27770
rect 14700 27718 14712 27770
rect 14712 27718 14742 27770
rect 14766 27718 14776 27770
rect 14776 27718 14822 27770
rect 14526 27716 14582 27718
rect 14606 27716 14662 27718
rect 14686 27716 14742 27718
rect 14766 27716 14822 27718
rect 19954 27770 20010 27772
rect 20034 27770 20090 27772
rect 20114 27770 20170 27772
rect 20194 27770 20250 27772
rect 19954 27718 20000 27770
rect 20000 27718 20010 27770
rect 20034 27718 20064 27770
rect 20064 27718 20076 27770
rect 20076 27718 20090 27770
rect 20114 27718 20128 27770
rect 20128 27718 20140 27770
rect 20140 27718 20170 27770
rect 20194 27718 20204 27770
rect 20204 27718 20250 27770
rect 19954 27716 20010 27718
rect 20034 27716 20090 27718
rect 20114 27716 20170 27718
rect 20194 27716 20250 27718
rect 6384 27226 6440 27228
rect 6464 27226 6520 27228
rect 6544 27226 6600 27228
rect 6624 27226 6680 27228
rect 6384 27174 6430 27226
rect 6430 27174 6440 27226
rect 6464 27174 6494 27226
rect 6494 27174 6506 27226
rect 6506 27174 6520 27226
rect 6544 27174 6558 27226
rect 6558 27174 6570 27226
rect 6570 27174 6600 27226
rect 6624 27174 6634 27226
rect 6634 27174 6680 27226
rect 6384 27172 6440 27174
rect 6464 27172 6520 27174
rect 6544 27172 6600 27174
rect 6624 27172 6680 27174
rect 11812 27226 11868 27228
rect 11892 27226 11948 27228
rect 11972 27226 12028 27228
rect 12052 27226 12108 27228
rect 11812 27174 11858 27226
rect 11858 27174 11868 27226
rect 11892 27174 11922 27226
rect 11922 27174 11934 27226
rect 11934 27174 11948 27226
rect 11972 27174 11986 27226
rect 11986 27174 11998 27226
rect 11998 27174 12028 27226
rect 12052 27174 12062 27226
rect 12062 27174 12108 27226
rect 11812 27172 11868 27174
rect 11892 27172 11948 27174
rect 11972 27172 12028 27174
rect 12052 27172 12108 27174
rect 17240 27226 17296 27228
rect 17320 27226 17376 27228
rect 17400 27226 17456 27228
rect 17480 27226 17536 27228
rect 17240 27174 17286 27226
rect 17286 27174 17296 27226
rect 17320 27174 17350 27226
rect 17350 27174 17362 27226
rect 17362 27174 17376 27226
rect 17400 27174 17414 27226
rect 17414 27174 17426 27226
rect 17426 27174 17456 27226
rect 17480 27174 17490 27226
rect 17490 27174 17536 27226
rect 17240 27172 17296 27174
rect 17320 27172 17376 27174
rect 17400 27172 17456 27174
rect 17480 27172 17536 27174
rect 22668 27226 22724 27228
rect 22748 27226 22804 27228
rect 22828 27226 22884 27228
rect 22908 27226 22964 27228
rect 22668 27174 22714 27226
rect 22714 27174 22724 27226
rect 22748 27174 22778 27226
rect 22778 27174 22790 27226
rect 22790 27174 22804 27226
rect 22828 27174 22842 27226
rect 22842 27174 22854 27226
rect 22854 27174 22884 27226
rect 22908 27174 22918 27226
rect 22918 27174 22964 27226
rect 22668 27172 22724 27174
rect 22748 27172 22804 27174
rect 22828 27172 22884 27174
rect 22908 27172 22964 27174
rect 22282 26852 22338 26888
rect 22282 26832 22284 26852
rect 22284 26832 22336 26852
rect 22336 26832 22338 26852
rect 3670 26682 3726 26684
rect 3750 26682 3806 26684
rect 3830 26682 3886 26684
rect 3910 26682 3966 26684
rect 3670 26630 3716 26682
rect 3716 26630 3726 26682
rect 3750 26630 3780 26682
rect 3780 26630 3792 26682
rect 3792 26630 3806 26682
rect 3830 26630 3844 26682
rect 3844 26630 3856 26682
rect 3856 26630 3886 26682
rect 3910 26630 3920 26682
rect 3920 26630 3966 26682
rect 3670 26628 3726 26630
rect 3750 26628 3806 26630
rect 3830 26628 3886 26630
rect 3910 26628 3966 26630
rect 9098 26682 9154 26684
rect 9178 26682 9234 26684
rect 9258 26682 9314 26684
rect 9338 26682 9394 26684
rect 9098 26630 9144 26682
rect 9144 26630 9154 26682
rect 9178 26630 9208 26682
rect 9208 26630 9220 26682
rect 9220 26630 9234 26682
rect 9258 26630 9272 26682
rect 9272 26630 9284 26682
rect 9284 26630 9314 26682
rect 9338 26630 9348 26682
rect 9348 26630 9394 26682
rect 9098 26628 9154 26630
rect 9178 26628 9234 26630
rect 9258 26628 9314 26630
rect 9338 26628 9394 26630
rect 14526 26682 14582 26684
rect 14606 26682 14662 26684
rect 14686 26682 14742 26684
rect 14766 26682 14822 26684
rect 14526 26630 14572 26682
rect 14572 26630 14582 26682
rect 14606 26630 14636 26682
rect 14636 26630 14648 26682
rect 14648 26630 14662 26682
rect 14686 26630 14700 26682
rect 14700 26630 14712 26682
rect 14712 26630 14742 26682
rect 14766 26630 14776 26682
rect 14776 26630 14822 26682
rect 14526 26628 14582 26630
rect 14606 26628 14662 26630
rect 14686 26628 14742 26630
rect 14766 26628 14822 26630
rect 19954 26682 20010 26684
rect 20034 26682 20090 26684
rect 20114 26682 20170 26684
rect 20194 26682 20250 26684
rect 19954 26630 20000 26682
rect 20000 26630 20010 26682
rect 20034 26630 20064 26682
rect 20064 26630 20076 26682
rect 20076 26630 20090 26682
rect 20114 26630 20128 26682
rect 20128 26630 20140 26682
rect 20140 26630 20170 26682
rect 20194 26630 20204 26682
rect 20204 26630 20250 26682
rect 19954 26628 20010 26630
rect 20034 26628 20090 26630
rect 20114 26628 20170 26630
rect 20194 26628 20250 26630
rect 22282 26324 22284 26344
rect 22284 26324 22336 26344
rect 22336 26324 22338 26344
rect 22282 26288 22338 26324
rect 1582 26152 1638 26208
rect 6384 26138 6440 26140
rect 6464 26138 6520 26140
rect 6544 26138 6600 26140
rect 6624 26138 6680 26140
rect 6384 26086 6430 26138
rect 6430 26086 6440 26138
rect 6464 26086 6494 26138
rect 6494 26086 6506 26138
rect 6506 26086 6520 26138
rect 6544 26086 6558 26138
rect 6558 26086 6570 26138
rect 6570 26086 6600 26138
rect 6624 26086 6634 26138
rect 6634 26086 6680 26138
rect 6384 26084 6440 26086
rect 6464 26084 6520 26086
rect 6544 26084 6600 26086
rect 6624 26084 6680 26086
rect 11812 26138 11868 26140
rect 11892 26138 11948 26140
rect 11972 26138 12028 26140
rect 12052 26138 12108 26140
rect 11812 26086 11858 26138
rect 11858 26086 11868 26138
rect 11892 26086 11922 26138
rect 11922 26086 11934 26138
rect 11934 26086 11948 26138
rect 11972 26086 11986 26138
rect 11986 26086 11998 26138
rect 11998 26086 12028 26138
rect 12052 26086 12062 26138
rect 12062 26086 12108 26138
rect 11812 26084 11868 26086
rect 11892 26084 11948 26086
rect 11972 26084 12028 26086
rect 12052 26084 12108 26086
rect 17240 26138 17296 26140
rect 17320 26138 17376 26140
rect 17400 26138 17456 26140
rect 17480 26138 17536 26140
rect 17240 26086 17286 26138
rect 17286 26086 17296 26138
rect 17320 26086 17350 26138
rect 17350 26086 17362 26138
rect 17362 26086 17376 26138
rect 17400 26086 17414 26138
rect 17414 26086 17426 26138
rect 17426 26086 17456 26138
rect 17480 26086 17490 26138
rect 17490 26086 17536 26138
rect 17240 26084 17296 26086
rect 17320 26084 17376 26086
rect 17400 26084 17456 26086
rect 17480 26084 17536 26086
rect 22668 26138 22724 26140
rect 22748 26138 22804 26140
rect 22828 26138 22884 26140
rect 22908 26138 22964 26140
rect 22668 26086 22714 26138
rect 22714 26086 22724 26138
rect 22748 26086 22778 26138
rect 22778 26086 22790 26138
rect 22790 26086 22804 26138
rect 22828 26086 22842 26138
rect 22842 26086 22854 26138
rect 22854 26086 22884 26138
rect 22908 26086 22918 26138
rect 22918 26086 22964 26138
rect 22668 26084 22724 26086
rect 22748 26084 22804 26086
rect 22828 26084 22884 26086
rect 22908 26084 22964 26086
rect 3670 25594 3726 25596
rect 3750 25594 3806 25596
rect 3830 25594 3886 25596
rect 3910 25594 3966 25596
rect 3670 25542 3716 25594
rect 3716 25542 3726 25594
rect 3750 25542 3780 25594
rect 3780 25542 3792 25594
rect 3792 25542 3806 25594
rect 3830 25542 3844 25594
rect 3844 25542 3856 25594
rect 3856 25542 3886 25594
rect 3910 25542 3920 25594
rect 3920 25542 3966 25594
rect 3670 25540 3726 25542
rect 3750 25540 3806 25542
rect 3830 25540 3886 25542
rect 3910 25540 3966 25542
rect 9098 25594 9154 25596
rect 9178 25594 9234 25596
rect 9258 25594 9314 25596
rect 9338 25594 9394 25596
rect 9098 25542 9144 25594
rect 9144 25542 9154 25594
rect 9178 25542 9208 25594
rect 9208 25542 9220 25594
rect 9220 25542 9234 25594
rect 9258 25542 9272 25594
rect 9272 25542 9284 25594
rect 9284 25542 9314 25594
rect 9338 25542 9348 25594
rect 9348 25542 9394 25594
rect 9098 25540 9154 25542
rect 9178 25540 9234 25542
rect 9258 25540 9314 25542
rect 9338 25540 9394 25542
rect 14526 25594 14582 25596
rect 14606 25594 14662 25596
rect 14686 25594 14742 25596
rect 14766 25594 14822 25596
rect 14526 25542 14572 25594
rect 14572 25542 14582 25594
rect 14606 25542 14636 25594
rect 14636 25542 14648 25594
rect 14648 25542 14662 25594
rect 14686 25542 14700 25594
rect 14700 25542 14712 25594
rect 14712 25542 14742 25594
rect 14766 25542 14776 25594
rect 14776 25542 14822 25594
rect 14526 25540 14582 25542
rect 14606 25540 14662 25542
rect 14686 25540 14742 25542
rect 14766 25540 14822 25542
rect 19954 25594 20010 25596
rect 20034 25594 20090 25596
rect 20114 25594 20170 25596
rect 20194 25594 20250 25596
rect 19954 25542 20000 25594
rect 20000 25542 20010 25594
rect 20034 25542 20064 25594
rect 20064 25542 20076 25594
rect 20076 25542 20090 25594
rect 20114 25542 20128 25594
rect 20128 25542 20140 25594
rect 20140 25542 20170 25594
rect 20194 25542 20204 25594
rect 20204 25542 20250 25594
rect 19954 25540 20010 25542
rect 20034 25540 20090 25542
rect 20114 25540 20170 25542
rect 20194 25540 20250 25542
rect 1582 25472 1638 25528
rect 22282 25236 22284 25256
rect 22284 25236 22336 25256
rect 22336 25236 22338 25256
rect 22282 25200 22338 25236
rect 6384 25050 6440 25052
rect 6464 25050 6520 25052
rect 6544 25050 6600 25052
rect 6624 25050 6680 25052
rect 6384 24998 6430 25050
rect 6430 24998 6440 25050
rect 6464 24998 6494 25050
rect 6494 24998 6506 25050
rect 6506 24998 6520 25050
rect 6544 24998 6558 25050
rect 6558 24998 6570 25050
rect 6570 24998 6600 25050
rect 6624 24998 6634 25050
rect 6634 24998 6680 25050
rect 6384 24996 6440 24998
rect 6464 24996 6520 24998
rect 6544 24996 6600 24998
rect 6624 24996 6680 24998
rect 11812 25050 11868 25052
rect 11892 25050 11948 25052
rect 11972 25050 12028 25052
rect 12052 25050 12108 25052
rect 11812 24998 11858 25050
rect 11858 24998 11868 25050
rect 11892 24998 11922 25050
rect 11922 24998 11934 25050
rect 11934 24998 11948 25050
rect 11972 24998 11986 25050
rect 11986 24998 11998 25050
rect 11998 24998 12028 25050
rect 12052 24998 12062 25050
rect 12062 24998 12108 25050
rect 11812 24996 11868 24998
rect 11892 24996 11948 24998
rect 11972 24996 12028 24998
rect 12052 24996 12108 24998
rect 17240 25050 17296 25052
rect 17320 25050 17376 25052
rect 17400 25050 17456 25052
rect 17480 25050 17536 25052
rect 17240 24998 17286 25050
rect 17286 24998 17296 25050
rect 17320 24998 17350 25050
rect 17350 24998 17362 25050
rect 17362 24998 17376 25050
rect 17400 24998 17414 25050
rect 17414 24998 17426 25050
rect 17426 24998 17456 25050
rect 17480 24998 17490 25050
rect 17490 24998 17536 25050
rect 17240 24996 17296 24998
rect 17320 24996 17376 24998
rect 17400 24996 17456 24998
rect 17480 24996 17536 24998
rect 22668 25050 22724 25052
rect 22748 25050 22804 25052
rect 22828 25050 22884 25052
rect 22908 25050 22964 25052
rect 22668 24998 22714 25050
rect 22714 24998 22724 25050
rect 22748 24998 22778 25050
rect 22778 24998 22790 25050
rect 22790 24998 22804 25050
rect 22828 24998 22842 25050
rect 22842 24998 22854 25050
rect 22854 24998 22884 25050
rect 22908 24998 22918 25050
rect 22918 24998 22964 25050
rect 22668 24996 22724 24998
rect 22748 24996 22804 24998
rect 22828 24996 22884 24998
rect 22908 24996 22964 24998
rect 22282 24676 22338 24712
rect 22282 24656 22284 24676
rect 22284 24656 22336 24676
rect 22336 24656 22338 24676
rect 3670 24506 3726 24508
rect 3750 24506 3806 24508
rect 3830 24506 3886 24508
rect 3910 24506 3966 24508
rect 3670 24454 3716 24506
rect 3716 24454 3726 24506
rect 3750 24454 3780 24506
rect 3780 24454 3792 24506
rect 3792 24454 3806 24506
rect 3830 24454 3844 24506
rect 3844 24454 3856 24506
rect 3856 24454 3886 24506
rect 3910 24454 3920 24506
rect 3920 24454 3966 24506
rect 3670 24452 3726 24454
rect 3750 24452 3806 24454
rect 3830 24452 3886 24454
rect 3910 24452 3966 24454
rect 9098 24506 9154 24508
rect 9178 24506 9234 24508
rect 9258 24506 9314 24508
rect 9338 24506 9394 24508
rect 9098 24454 9144 24506
rect 9144 24454 9154 24506
rect 9178 24454 9208 24506
rect 9208 24454 9220 24506
rect 9220 24454 9234 24506
rect 9258 24454 9272 24506
rect 9272 24454 9284 24506
rect 9284 24454 9314 24506
rect 9338 24454 9348 24506
rect 9348 24454 9394 24506
rect 9098 24452 9154 24454
rect 9178 24452 9234 24454
rect 9258 24452 9314 24454
rect 9338 24452 9394 24454
rect 14526 24506 14582 24508
rect 14606 24506 14662 24508
rect 14686 24506 14742 24508
rect 14766 24506 14822 24508
rect 14526 24454 14572 24506
rect 14572 24454 14582 24506
rect 14606 24454 14636 24506
rect 14636 24454 14648 24506
rect 14648 24454 14662 24506
rect 14686 24454 14700 24506
rect 14700 24454 14712 24506
rect 14712 24454 14742 24506
rect 14766 24454 14776 24506
rect 14776 24454 14822 24506
rect 14526 24452 14582 24454
rect 14606 24452 14662 24454
rect 14686 24452 14742 24454
rect 14766 24452 14822 24454
rect 19954 24506 20010 24508
rect 20034 24506 20090 24508
rect 20114 24506 20170 24508
rect 20194 24506 20250 24508
rect 19954 24454 20000 24506
rect 20000 24454 20010 24506
rect 20034 24454 20064 24506
rect 20064 24454 20076 24506
rect 20076 24454 20090 24506
rect 20114 24454 20128 24506
rect 20128 24454 20140 24506
rect 20140 24454 20170 24506
rect 20194 24454 20204 24506
rect 20204 24454 20250 24506
rect 19954 24452 20010 24454
rect 20034 24452 20090 24454
rect 20114 24452 20170 24454
rect 20194 24452 20250 24454
rect 1582 24148 1584 24168
rect 1584 24148 1636 24168
rect 1636 24148 1638 24168
rect 1582 24112 1638 24148
rect 6384 23962 6440 23964
rect 6464 23962 6520 23964
rect 6544 23962 6600 23964
rect 6624 23962 6680 23964
rect 6384 23910 6430 23962
rect 6430 23910 6440 23962
rect 6464 23910 6494 23962
rect 6494 23910 6506 23962
rect 6506 23910 6520 23962
rect 6544 23910 6558 23962
rect 6558 23910 6570 23962
rect 6570 23910 6600 23962
rect 6624 23910 6634 23962
rect 6634 23910 6680 23962
rect 6384 23908 6440 23910
rect 6464 23908 6520 23910
rect 6544 23908 6600 23910
rect 6624 23908 6680 23910
rect 11812 23962 11868 23964
rect 11892 23962 11948 23964
rect 11972 23962 12028 23964
rect 12052 23962 12108 23964
rect 11812 23910 11858 23962
rect 11858 23910 11868 23962
rect 11892 23910 11922 23962
rect 11922 23910 11934 23962
rect 11934 23910 11948 23962
rect 11972 23910 11986 23962
rect 11986 23910 11998 23962
rect 11998 23910 12028 23962
rect 12052 23910 12062 23962
rect 12062 23910 12108 23962
rect 11812 23908 11868 23910
rect 11892 23908 11948 23910
rect 11972 23908 12028 23910
rect 12052 23908 12108 23910
rect 17240 23962 17296 23964
rect 17320 23962 17376 23964
rect 17400 23962 17456 23964
rect 17480 23962 17536 23964
rect 17240 23910 17286 23962
rect 17286 23910 17296 23962
rect 17320 23910 17350 23962
rect 17350 23910 17362 23962
rect 17362 23910 17376 23962
rect 17400 23910 17414 23962
rect 17414 23910 17426 23962
rect 17426 23910 17456 23962
rect 17480 23910 17490 23962
rect 17490 23910 17536 23962
rect 17240 23908 17296 23910
rect 17320 23908 17376 23910
rect 17400 23908 17456 23910
rect 17480 23908 17536 23910
rect 22668 23962 22724 23964
rect 22748 23962 22804 23964
rect 22828 23962 22884 23964
rect 22908 23962 22964 23964
rect 22668 23910 22714 23962
rect 22714 23910 22724 23962
rect 22748 23910 22778 23962
rect 22778 23910 22790 23962
rect 22790 23910 22804 23962
rect 22828 23910 22842 23962
rect 22842 23910 22854 23962
rect 22854 23910 22884 23962
rect 22908 23910 22918 23962
rect 22918 23910 22964 23962
rect 22668 23908 22724 23910
rect 22748 23908 22804 23910
rect 22828 23908 22884 23910
rect 22908 23908 22964 23910
rect 22282 23588 22338 23624
rect 22282 23568 22284 23588
rect 22284 23568 22336 23588
rect 22336 23568 22338 23588
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 3670 23418 3726 23420
rect 3750 23418 3806 23420
rect 3830 23418 3886 23420
rect 3910 23418 3966 23420
rect 3670 23366 3716 23418
rect 3716 23366 3726 23418
rect 3750 23366 3780 23418
rect 3780 23366 3792 23418
rect 3792 23366 3806 23418
rect 3830 23366 3844 23418
rect 3844 23366 3856 23418
rect 3856 23366 3886 23418
rect 3910 23366 3920 23418
rect 3920 23366 3966 23418
rect 3670 23364 3726 23366
rect 3750 23364 3806 23366
rect 3830 23364 3886 23366
rect 3910 23364 3966 23366
rect 9098 23418 9154 23420
rect 9178 23418 9234 23420
rect 9258 23418 9314 23420
rect 9338 23418 9394 23420
rect 9098 23366 9144 23418
rect 9144 23366 9154 23418
rect 9178 23366 9208 23418
rect 9208 23366 9220 23418
rect 9220 23366 9234 23418
rect 9258 23366 9272 23418
rect 9272 23366 9284 23418
rect 9284 23366 9314 23418
rect 9338 23366 9348 23418
rect 9348 23366 9394 23418
rect 9098 23364 9154 23366
rect 9178 23364 9234 23366
rect 9258 23364 9314 23366
rect 9338 23364 9394 23366
rect 14526 23418 14582 23420
rect 14606 23418 14662 23420
rect 14686 23418 14742 23420
rect 14766 23418 14822 23420
rect 14526 23366 14572 23418
rect 14572 23366 14582 23418
rect 14606 23366 14636 23418
rect 14636 23366 14648 23418
rect 14648 23366 14662 23418
rect 14686 23366 14700 23418
rect 14700 23366 14712 23418
rect 14712 23366 14742 23418
rect 14766 23366 14776 23418
rect 14776 23366 14822 23418
rect 14526 23364 14582 23366
rect 14606 23364 14662 23366
rect 14686 23364 14742 23366
rect 14766 23364 14822 23366
rect 19954 23418 20010 23420
rect 20034 23418 20090 23420
rect 20114 23418 20170 23420
rect 20194 23418 20250 23420
rect 19954 23366 20000 23418
rect 20000 23366 20010 23418
rect 20034 23366 20064 23418
rect 20064 23366 20076 23418
rect 20076 23366 20090 23418
rect 20114 23366 20128 23418
rect 20128 23366 20140 23418
rect 20140 23366 20170 23418
rect 20194 23366 20204 23418
rect 20204 23366 20250 23418
rect 19954 23364 20010 23366
rect 20034 23364 20090 23366
rect 20114 23364 20170 23366
rect 20194 23364 20250 23366
rect 22282 23060 22284 23080
rect 22284 23060 22336 23080
rect 22336 23060 22338 23080
rect 22282 23024 22338 23060
rect 6384 22874 6440 22876
rect 6464 22874 6520 22876
rect 6544 22874 6600 22876
rect 6624 22874 6680 22876
rect 6384 22822 6430 22874
rect 6430 22822 6440 22874
rect 6464 22822 6494 22874
rect 6494 22822 6506 22874
rect 6506 22822 6520 22874
rect 6544 22822 6558 22874
rect 6558 22822 6570 22874
rect 6570 22822 6600 22874
rect 6624 22822 6634 22874
rect 6634 22822 6680 22874
rect 6384 22820 6440 22822
rect 6464 22820 6520 22822
rect 6544 22820 6600 22822
rect 6624 22820 6680 22822
rect 11812 22874 11868 22876
rect 11892 22874 11948 22876
rect 11972 22874 12028 22876
rect 12052 22874 12108 22876
rect 11812 22822 11858 22874
rect 11858 22822 11868 22874
rect 11892 22822 11922 22874
rect 11922 22822 11934 22874
rect 11934 22822 11948 22874
rect 11972 22822 11986 22874
rect 11986 22822 11998 22874
rect 11998 22822 12028 22874
rect 12052 22822 12062 22874
rect 12062 22822 12108 22874
rect 11812 22820 11868 22822
rect 11892 22820 11948 22822
rect 11972 22820 12028 22822
rect 12052 22820 12108 22822
rect 17240 22874 17296 22876
rect 17320 22874 17376 22876
rect 17400 22874 17456 22876
rect 17480 22874 17536 22876
rect 17240 22822 17286 22874
rect 17286 22822 17296 22874
rect 17320 22822 17350 22874
rect 17350 22822 17362 22874
rect 17362 22822 17376 22874
rect 17400 22822 17414 22874
rect 17414 22822 17426 22874
rect 17426 22822 17456 22874
rect 17480 22822 17490 22874
rect 17490 22822 17536 22874
rect 17240 22820 17296 22822
rect 17320 22820 17376 22822
rect 17400 22820 17456 22822
rect 17480 22820 17536 22822
rect 22668 22874 22724 22876
rect 22748 22874 22804 22876
rect 22828 22874 22884 22876
rect 22908 22874 22964 22876
rect 22668 22822 22714 22874
rect 22714 22822 22724 22874
rect 22748 22822 22778 22874
rect 22778 22822 22790 22874
rect 22790 22822 22804 22874
rect 22828 22822 22842 22874
rect 22842 22822 22854 22874
rect 22854 22822 22884 22874
rect 22908 22822 22918 22874
rect 22918 22822 22964 22874
rect 22668 22820 22724 22822
rect 22748 22820 22804 22822
rect 22828 22820 22884 22822
rect 22908 22820 22964 22822
rect 3670 22330 3726 22332
rect 3750 22330 3806 22332
rect 3830 22330 3886 22332
rect 3910 22330 3966 22332
rect 3670 22278 3716 22330
rect 3716 22278 3726 22330
rect 3750 22278 3780 22330
rect 3780 22278 3792 22330
rect 3792 22278 3806 22330
rect 3830 22278 3844 22330
rect 3844 22278 3856 22330
rect 3856 22278 3886 22330
rect 3910 22278 3920 22330
rect 3920 22278 3966 22330
rect 3670 22276 3726 22278
rect 3750 22276 3806 22278
rect 3830 22276 3886 22278
rect 3910 22276 3966 22278
rect 9098 22330 9154 22332
rect 9178 22330 9234 22332
rect 9258 22330 9314 22332
rect 9338 22330 9394 22332
rect 9098 22278 9144 22330
rect 9144 22278 9154 22330
rect 9178 22278 9208 22330
rect 9208 22278 9220 22330
rect 9220 22278 9234 22330
rect 9258 22278 9272 22330
rect 9272 22278 9284 22330
rect 9284 22278 9314 22330
rect 9338 22278 9348 22330
rect 9348 22278 9394 22330
rect 9098 22276 9154 22278
rect 9178 22276 9234 22278
rect 9258 22276 9314 22278
rect 9338 22276 9394 22278
rect 14526 22330 14582 22332
rect 14606 22330 14662 22332
rect 14686 22330 14742 22332
rect 14766 22330 14822 22332
rect 14526 22278 14572 22330
rect 14572 22278 14582 22330
rect 14606 22278 14636 22330
rect 14636 22278 14648 22330
rect 14648 22278 14662 22330
rect 14686 22278 14700 22330
rect 14700 22278 14712 22330
rect 14712 22278 14742 22330
rect 14766 22278 14776 22330
rect 14776 22278 14822 22330
rect 14526 22276 14582 22278
rect 14606 22276 14662 22278
rect 14686 22276 14742 22278
rect 14766 22276 14822 22278
rect 19954 22330 20010 22332
rect 20034 22330 20090 22332
rect 20114 22330 20170 22332
rect 20194 22330 20250 22332
rect 19954 22278 20000 22330
rect 20000 22278 20010 22330
rect 20034 22278 20064 22330
rect 20064 22278 20076 22330
rect 20076 22278 20090 22330
rect 20114 22278 20128 22330
rect 20128 22278 20140 22330
rect 20140 22278 20170 22330
rect 20194 22278 20204 22330
rect 20204 22278 20250 22330
rect 19954 22276 20010 22278
rect 20034 22276 20090 22278
rect 20114 22276 20170 22278
rect 20194 22276 20250 22278
rect 1582 22072 1638 22128
rect 22282 21936 22338 21992
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 1582 21428 1584 21448
rect 1584 21428 1636 21448
rect 1636 21428 1638 21448
rect 1582 21392 1638 21428
rect 22282 21412 22338 21448
rect 22282 21392 22284 21412
rect 22284 21392 22336 21412
rect 22336 21392 22338 21412
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 22282 20324 22338 20360
rect 22282 20304 22284 20324
rect 22284 20304 22336 20324
rect 22336 20304 22338 20324
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 1582 20032 1638 20088
rect 22282 19796 22284 19816
rect 22284 19796 22336 19816
rect 22336 19796 22338 19816
rect 22282 19760 22338 19796
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 1582 19352 1638 19408
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 22282 18708 22284 18728
rect 22284 18708 22336 18728
rect 22336 18708 22338 18728
rect 22282 18672 22338 18708
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 22282 18148 22338 18184
rect 22282 18128 22284 18148
rect 22284 18128 22336 18148
rect 22336 18128 22338 18148
rect 1582 18028 1584 18048
rect 1584 18028 1636 18048
rect 1636 18028 1638 18048
rect 1582 17992 1638 18028
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 1582 17312 1638 17368
rect 22282 17060 22338 17096
rect 22282 17040 22284 17060
rect 22284 17040 22336 17060
rect 22336 17040 22338 17060
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 22282 16496 22338 16552
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 1582 15988 1584 16008
rect 1584 15988 1636 16008
rect 1636 15988 1638 16008
rect 1582 15952 1638 15988
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 22282 15444 22284 15464
rect 22284 15444 22336 15464
rect 22336 15444 22338 15464
rect 22282 15408 22338 15444
rect 1582 15272 1638 15328
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 22282 14884 22338 14920
rect 22282 14864 22284 14884
rect 22284 14864 22336 14884
rect 22336 14864 22338 14884
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 1582 13912 1638 13968
rect 22282 13812 22284 13832
rect 22284 13812 22336 13832
rect 22336 13812 22338 13832
rect 22282 13776 22338 13812
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 1582 13268 1584 13288
rect 1584 13268 1636 13288
rect 1636 13268 1638 13288
rect 1582 13232 1638 13268
rect 22282 13268 22284 13288
rect 22284 13268 22336 13288
rect 22336 13268 22338 13288
rect 22282 13232 22338 13268
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 22282 12180 22284 12200
rect 22284 12180 22336 12200
rect 22336 12180 22338 12200
rect 22282 12144 22338 12180
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 1582 11872 1638 11928
rect 22282 11620 22338 11656
rect 22282 11600 22284 11620
rect 22284 11600 22336 11620
rect 22336 11600 22338 11620
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 1582 11192 1638 11248
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 22282 10532 22338 10568
rect 22282 10512 22284 10532
rect 22284 10512 22336 10532
rect 22336 10512 22338 10532
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 22282 10004 22284 10024
rect 22284 10004 22336 10024
rect 22336 10004 22338 10024
rect 22282 9968 22338 10004
rect 1582 9832 1638 9888
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 1582 9152 1638 9208
rect 22282 8916 22284 8936
rect 22284 8916 22336 8936
rect 22336 8916 22338 8936
rect 22282 8880 22338 8916
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 22282 8356 22338 8392
rect 22282 8336 22284 8356
rect 22284 8336 22336 8356
rect 22336 8336 22338 8356
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 1582 7828 1584 7848
rect 1584 7828 1636 7848
rect 1636 7828 1638 7848
rect 1582 7792 1638 7828
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 22282 7268 22338 7304
rect 22282 7248 22284 7268
rect 22284 7248 22336 7268
rect 22336 7248 22338 7268
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 22282 6740 22284 6760
rect 22284 6740 22336 6760
rect 22336 6740 22338 6760
rect 22282 6704 22338 6740
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 1582 5752 1638 5808
rect 22282 5652 22284 5672
rect 22284 5652 22336 5672
rect 22336 5652 22338 5672
rect 22282 5616 22338 5652
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 1582 5108 1584 5128
rect 1584 5108 1636 5128
rect 1636 5108 1638 5128
rect 1582 5072 1638 5108
rect 22282 5092 22338 5128
rect 22282 5072 22284 5092
rect 22284 5072 22336 5092
rect 22336 5072 22338 5092
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 22282 4004 22338 4040
rect 22282 3984 22284 4004
rect 22284 3984 22336 4004
rect 22336 3984 22338 4004
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 1582 3712 1638 3768
rect 22282 3476 22284 3496
rect 22284 3476 22336 3496
rect 22336 3476 22338 3496
rect 22282 3440 22338 3476
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 1582 3032 1638 3088
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
rect 1582 1672 1638 1728
rect 1398 992 1454 1048
<< metal3 >>
rect 0 28840 800 28960
rect 0 28250 800 28280
rect 2865 28250 2931 28253
rect 0 28248 2931 28250
rect 0 28192 2870 28248
rect 2926 28192 2931 28248
rect 0 28190 2931 28192
rect 0 28160 800 28190
rect 2865 28187 2931 28190
rect 3660 27776 3976 27777
rect 3660 27712 3666 27776
rect 3730 27712 3746 27776
rect 3810 27712 3826 27776
rect 3890 27712 3906 27776
rect 3970 27712 3976 27776
rect 3660 27711 3976 27712
rect 9088 27776 9404 27777
rect 9088 27712 9094 27776
rect 9158 27712 9174 27776
rect 9238 27712 9254 27776
rect 9318 27712 9334 27776
rect 9398 27712 9404 27776
rect 9088 27711 9404 27712
rect 14516 27776 14832 27777
rect 14516 27712 14522 27776
rect 14586 27712 14602 27776
rect 14666 27712 14682 27776
rect 14746 27712 14762 27776
rect 14826 27712 14832 27776
rect 14516 27711 14832 27712
rect 19944 27776 20260 27777
rect 19944 27712 19950 27776
rect 20014 27712 20030 27776
rect 20094 27712 20110 27776
rect 20174 27712 20190 27776
rect 20254 27712 20260 27776
rect 19944 27711 20260 27712
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 6374 27232 6690 27233
rect 6374 27168 6380 27232
rect 6444 27168 6460 27232
rect 6524 27168 6540 27232
rect 6604 27168 6620 27232
rect 6684 27168 6690 27232
rect 6374 27167 6690 27168
rect 11802 27232 12118 27233
rect 11802 27168 11808 27232
rect 11872 27168 11888 27232
rect 11952 27168 11968 27232
rect 12032 27168 12048 27232
rect 12112 27168 12118 27232
rect 11802 27167 12118 27168
rect 17230 27232 17546 27233
rect 17230 27168 17236 27232
rect 17300 27168 17316 27232
rect 17380 27168 17396 27232
rect 17460 27168 17476 27232
rect 17540 27168 17546 27232
rect 17230 27167 17546 27168
rect 22658 27232 22974 27233
rect 22658 27168 22664 27232
rect 22728 27168 22744 27232
rect 22808 27168 22824 27232
rect 22888 27168 22904 27232
rect 22968 27168 22974 27232
rect 22658 27167 22974 27168
rect 0 26800 800 26920
rect 22277 26890 22343 26893
rect 23200 26890 24000 26920
rect 22277 26888 24000 26890
rect 22277 26832 22282 26888
rect 22338 26832 24000 26888
rect 22277 26830 24000 26832
rect 22277 26827 22343 26830
rect 23200 26800 24000 26830
rect 3660 26688 3976 26689
rect 3660 26624 3666 26688
rect 3730 26624 3746 26688
rect 3810 26624 3826 26688
rect 3890 26624 3906 26688
rect 3970 26624 3976 26688
rect 3660 26623 3976 26624
rect 9088 26688 9404 26689
rect 9088 26624 9094 26688
rect 9158 26624 9174 26688
rect 9238 26624 9254 26688
rect 9318 26624 9334 26688
rect 9398 26624 9404 26688
rect 9088 26623 9404 26624
rect 14516 26688 14832 26689
rect 14516 26624 14522 26688
rect 14586 26624 14602 26688
rect 14666 26624 14682 26688
rect 14746 26624 14762 26688
rect 14826 26624 14832 26688
rect 14516 26623 14832 26624
rect 19944 26688 20260 26689
rect 19944 26624 19950 26688
rect 20014 26624 20030 26688
rect 20094 26624 20110 26688
rect 20174 26624 20190 26688
rect 20254 26624 20260 26688
rect 19944 26623 20260 26624
rect 22277 26346 22343 26349
rect 23200 26346 24000 26376
rect 22277 26344 24000 26346
rect 22277 26288 22282 26344
rect 22338 26288 24000 26344
rect 22277 26286 24000 26288
rect 22277 26283 22343 26286
rect 23200 26256 24000 26286
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 6374 26144 6690 26145
rect 6374 26080 6380 26144
rect 6444 26080 6460 26144
rect 6524 26080 6540 26144
rect 6604 26080 6620 26144
rect 6684 26080 6690 26144
rect 6374 26079 6690 26080
rect 11802 26144 12118 26145
rect 11802 26080 11808 26144
rect 11872 26080 11888 26144
rect 11952 26080 11968 26144
rect 12032 26080 12048 26144
rect 12112 26080 12118 26144
rect 11802 26079 12118 26080
rect 17230 26144 17546 26145
rect 17230 26080 17236 26144
rect 17300 26080 17316 26144
rect 17380 26080 17396 26144
rect 17460 26080 17476 26144
rect 17540 26080 17546 26144
rect 17230 26079 17546 26080
rect 22658 26144 22974 26145
rect 22658 26080 22664 26144
rect 22728 26080 22744 26144
rect 22808 26080 22824 26144
rect 22888 26080 22904 26144
rect 22968 26080 22974 26144
rect 22658 26079 22974 26080
rect 23200 25712 24000 25832
rect 3660 25600 3976 25601
rect 0 25530 800 25560
rect 3660 25536 3666 25600
rect 3730 25536 3746 25600
rect 3810 25536 3826 25600
rect 3890 25536 3906 25600
rect 3970 25536 3976 25600
rect 3660 25535 3976 25536
rect 9088 25600 9404 25601
rect 9088 25536 9094 25600
rect 9158 25536 9174 25600
rect 9238 25536 9254 25600
rect 9318 25536 9334 25600
rect 9398 25536 9404 25600
rect 9088 25535 9404 25536
rect 14516 25600 14832 25601
rect 14516 25536 14522 25600
rect 14586 25536 14602 25600
rect 14666 25536 14682 25600
rect 14746 25536 14762 25600
rect 14826 25536 14832 25600
rect 14516 25535 14832 25536
rect 19944 25600 20260 25601
rect 19944 25536 19950 25600
rect 20014 25536 20030 25600
rect 20094 25536 20110 25600
rect 20174 25536 20190 25600
rect 20254 25536 20260 25600
rect 19944 25535 20260 25536
rect 1577 25530 1643 25533
rect 0 25528 1643 25530
rect 0 25472 1582 25528
rect 1638 25472 1643 25528
rect 0 25470 1643 25472
rect 0 25440 800 25470
rect 1577 25467 1643 25470
rect 22277 25258 22343 25261
rect 23200 25258 24000 25288
rect 22277 25256 24000 25258
rect 22277 25200 22282 25256
rect 22338 25200 24000 25256
rect 22277 25198 24000 25200
rect 22277 25195 22343 25198
rect 23200 25168 24000 25198
rect 6374 25056 6690 25057
rect 6374 24992 6380 25056
rect 6444 24992 6460 25056
rect 6524 24992 6540 25056
rect 6604 24992 6620 25056
rect 6684 24992 6690 25056
rect 6374 24991 6690 24992
rect 11802 25056 12118 25057
rect 11802 24992 11808 25056
rect 11872 24992 11888 25056
rect 11952 24992 11968 25056
rect 12032 24992 12048 25056
rect 12112 24992 12118 25056
rect 11802 24991 12118 24992
rect 17230 25056 17546 25057
rect 17230 24992 17236 25056
rect 17300 24992 17316 25056
rect 17380 24992 17396 25056
rect 17460 24992 17476 25056
rect 17540 24992 17546 25056
rect 17230 24991 17546 24992
rect 22658 25056 22974 25057
rect 22658 24992 22664 25056
rect 22728 24992 22744 25056
rect 22808 24992 22824 25056
rect 22888 24992 22904 25056
rect 22968 24992 22974 25056
rect 22658 24991 22974 24992
rect 0 24760 800 24880
rect 22277 24714 22343 24717
rect 23200 24714 24000 24744
rect 22277 24712 24000 24714
rect 22277 24656 22282 24712
rect 22338 24656 24000 24712
rect 22277 24654 24000 24656
rect 22277 24651 22343 24654
rect 23200 24624 24000 24654
rect 3660 24512 3976 24513
rect 3660 24448 3666 24512
rect 3730 24448 3746 24512
rect 3810 24448 3826 24512
rect 3890 24448 3906 24512
rect 3970 24448 3976 24512
rect 3660 24447 3976 24448
rect 9088 24512 9404 24513
rect 9088 24448 9094 24512
rect 9158 24448 9174 24512
rect 9238 24448 9254 24512
rect 9318 24448 9334 24512
rect 9398 24448 9404 24512
rect 9088 24447 9404 24448
rect 14516 24512 14832 24513
rect 14516 24448 14522 24512
rect 14586 24448 14602 24512
rect 14666 24448 14682 24512
rect 14746 24448 14762 24512
rect 14826 24448 14832 24512
rect 14516 24447 14832 24448
rect 19944 24512 20260 24513
rect 19944 24448 19950 24512
rect 20014 24448 20030 24512
rect 20094 24448 20110 24512
rect 20174 24448 20190 24512
rect 20254 24448 20260 24512
rect 19944 24447 20260 24448
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 23200 24080 24000 24200
rect 6374 23968 6690 23969
rect 6374 23904 6380 23968
rect 6444 23904 6460 23968
rect 6524 23904 6540 23968
rect 6604 23904 6620 23968
rect 6684 23904 6690 23968
rect 6374 23903 6690 23904
rect 11802 23968 12118 23969
rect 11802 23904 11808 23968
rect 11872 23904 11888 23968
rect 11952 23904 11968 23968
rect 12032 23904 12048 23968
rect 12112 23904 12118 23968
rect 11802 23903 12118 23904
rect 17230 23968 17546 23969
rect 17230 23904 17236 23968
rect 17300 23904 17316 23968
rect 17380 23904 17396 23968
rect 17460 23904 17476 23968
rect 17540 23904 17546 23968
rect 17230 23903 17546 23904
rect 22658 23968 22974 23969
rect 22658 23904 22664 23968
rect 22728 23904 22744 23968
rect 22808 23904 22824 23968
rect 22888 23904 22904 23968
rect 22968 23904 22974 23968
rect 22658 23903 22974 23904
rect 22277 23626 22343 23629
rect 23200 23626 24000 23656
rect 22277 23624 24000 23626
rect 22277 23568 22282 23624
rect 22338 23568 24000 23624
rect 22277 23566 24000 23568
rect 22277 23563 22343 23566
rect 23200 23536 24000 23566
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 3660 23424 3976 23425
rect 3660 23360 3666 23424
rect 3730 23360 3746 23424
rect 3810 23360 3826 23424
rect 3890 23360 3906 23424
rect 3970 23360 3976 23424
rect 3660 23359 3976 23360
rect 9088 23424 9404 23425
rect 9088 23360 9094 23424
rect 9158 23360 9174 23424
rect 9238 23360 9254 23424
rect 9318 23360 9334 23424
rect 9398 23360 9404 23424
rect 9088 23359 9404 23360
rect 14516 23424 14832 23425
rect 14516 23360 14522 23424
rect 14586 23360 14602 23424
rect 14666 23360 14682 23424
rect 14746 23360 14762 23424
rect 14826 23360 14832 23424
rect 14516 23359 14832 23360
rect 19944 23424 20260 23425
rect 19944 23360 19950 23424
rect 20014 23360 20030 23424
rect 20094 23360 20110 23424
rect 20174 23360 20190 23424
rect 20254 23360 20260 23424
rect 19944 23359 20260 23360
rect 22277 23082 22343 23085
rect 23200 23082 24000 23112
rect 22277 23080 24000 23082
rect 22277 23024 22282 23080
rect 22338 23024 24000 23080
rect 22277 23022 24000 23024
rect 22277 23019 22343 23022
rect 23200 22992 24000 23022
rect 6374 22880 6690 22881
rect 0 22720 800 22840
rect 6374 22816 6380 22880
rect 6444 22816 6460 22880
rect 6524 22816 6540 22880
rect 6604 22816 6620 22880
rect 6684 22816 6690 22880
rect 6374 22815 6690 22816
rect 11802 22880 12118 22881
rect 11802 22816 11808 22880
rect 11872 22816 11888 22880
rect 11952 22816 11968 22880
rect 12032 22816 12048 22880
rect 12112 22816 12118 22880
rect 11802 22815 12118 22816
rect 17230 22880 17546 22881
rect 17230 22816 17236 22880
rect 17300 22816 17316 22880
rect 17380 22816 17396 22880
rect 17460 22816 17476 22880
rect 17540 22816 17546 22880
rect 17230 22815 17546 22816
rect 22658 22880 22974 22881
rect 22658 22816 22664 22880
rect 22728 22816 22744 22880
rect 22808 22816 22824 22880
rect 22888 22816 22904 22880
rect 22968 22816 22974 22880
rect 22658 22815 22974 22816
rect 23200 22448 24000 22568
rect 3660 22336 3976 22337
rect 3660 22272 3666 22336
rect 3730 22272 3746 22336
rect 3810 22272 3826 22336
rect 3890 22272 3906 22336
rect 3970 22272 3976 22336
rect 3660 22271 3976 22272
rect 9088 22336 9404 22337
rect 9088 22272 9094 22336
rect 9158 22272 9174 22336
rect 9238 22272 9254 22336
rect 9318 22272 9334 22336
rect 9398 22272 9404 22336
rect 9088 22271 9404 22272
rect 14516 22336 14832 22337
rect 14516 22272 14522 22336
rect 14586 22272 14602 22336
rect 14666 22272 14682 22336
rect 14746 22272 14762 22336
rect 14826 22272 14832 22336
rect 14516 22271 14832 22272
rect 19944 22336 20260 22337
rect 19944 22272 19950 22336
rect 20014 22272 20030 22336
rect 20094 22272 20110 22336
rect 20174 22272 20190 22336
rect 20254 22272 20260 22336
rect 19944 22271 20260 22272
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 22277 21994 22343 21997
rect 23200 21994 24000 22024
rect 22277 21992 24000 21994
rect 22277 21936 22282 21992
rect 22338 21936 24000 21992
rect 22277 21934 24000 21936
rect 22277 21931 22343 21934
rect 23200 21904 24000 21934
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 22277 21450 22343 21453
rect 23200 21450 24000 21480
rect 22277 21448 24000 21450
rect 22277 21392 22282 21448
rect 22338 21392 24000 21448
rect 22277 21390 24000 21392
rect 22277 21387 22343 21390
rect 23200 21360 24000 21390
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 23200 20816 24000 20936
rect 0 20680 800 20800
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 22277 20362 22343 20365
rect 23200 20362 24000 20392
rect 22277 20360 24000 20362
rect 22277 20304 22282 20360
rect 22338 20304 24000 20360
rect 22277 20302 24000 20304
rect 22277 20299 22343 20302
rect 23200 20272 24000 20302
rect 3660 20160 3976 20161
rect 0 20090 800 20120
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 22277 19818 22343 19821
rect 23200 19818 24000 19848
rect 22277 19816 24000 19818
rect 22277 19760 22282 19816
rect 22338 19760 24000 19816
rect 22277 19758 24000 19760
rect 22277 19755 22343 19758
rect 23200 19728 24000 19758
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 23200 19184 24000 19304
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 0 18640 800 18760
rect 22277 18730 22343 18733
rect 23200 18730 24000 18760
rect 22277 18728 24000 18730
rect 22277 18672 22282 18728
rect 22338 18672 24000 18728
rect 22277 18670 24000 18672
rect 22277 18667 22343 18670
rect 23200 18640 24000 18670
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 22277 18186 22343 18189
rect 23200 18186 24000 18216
rect 22277 18184 24000 18186
rect 22277 18128 22282 18184
rect 22338 18128 24000 18184
rect 22277 18126 24000 18128
rect 22277 18123 22343 18126
rect 23200 18096 24000 18126
rect 0 18050 800 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 800 17990
rect 1577 17987 1643 17990
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 23200 17552 24000 17672
rect 6374 17440 6690 17441
rect 0 17370 800 17400
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 22277 17098 22343 17101
rect 23200 17098 24000 17128
rect 22277 17096 24000 17098
rect 22277 17040 22282 17096
rect 22338 17040 24000 17096
rect 22277 17038 24000 17040
rect 22277 17035 22343 17038
rect 23200 17008 24000 17038
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 0 16600 800 16720
rect 22277 16554 22343 16557
rect 23200 16554 24000 16584
rect 22277 16552 24000 16554
rect 22277 16496 22282 16552
rect 22338 16496 24000 16552
rect 22277 16494 24000 16496
rect 22277 16491 22343 16494
rect 23200 16464 24000 16494
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 0 16010 800 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 800 15950
rect 1577 15947 1643 15950
rect 23200 15920 24000 16040
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 22277 15466 22343 15469
rect 23200 15466 24000 15496
rect 22277 15464 24000 15466
rect 22277 15408 22282 15464
rect 22338 15408 24000 15464
rect 22277 15406 24000 15408
rect 22277 15403 22343 15406
rect 23200 15376 24000 15406
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 22277 14922 22343 14925
rect 23200 14922 24000 14952
rect 22277 14920 24000 14922
rect 22277 14864 22282 14920
rect 22338 14864 24000 14920
rect 22277 14862 24000 14864
rect 22277 14859 22343 14862
rect 23200 14832 24000 14862
rect 3660 14720 3976 14721
rect 0 14560 800 14680
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 23200 14288 24000 14408
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 22277 13834 22343 13837
rect 23200 13834 24000 13864
rect 22277 13832 24000 13834
rect 22277 13776 22282 13832
rect 22338 13776 24000 13832
rect 22277 13774 24000 13776
rect 22277 13771 22343 13774
rect 23200 13744 24000 13774
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 22277 13290 22343 13293
rect 23200 13290 24000 13320
rect 22277 13288 24000 13290
rect 22277 13232 22282 13288
rect 22338 13232 24000 13288
rect 22277 13230 24000 13232
rect 22277 13227 22343 13230
rect 23200 13200 24000 13230
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 23200 12656 24000 12776
rect 0 12520 800 12640
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 22277 12202 22343 12205
rect 23200 12202 24000 12232
rect 22277 12200 24000 12202
rect 22277 12144 22282 12200
rect 22338 12144 24000 12200
rect 22277 12142 24000 12144
rect 22277 12139 22343 12142
rect 23200 12112 24000 12142
rect 6374 12000 6690 12001
rect 0 11930 800 11960
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 800 11870
rect 1577 11867 1643 11870
rect 22277 11658 22343 11661
rect 23200 11658 24000 11688
rect 22277 11656 24000 11658
rect 22277 11600 22282 11656
rect 22338 11600 24000 11656
rect 22277 11598 24000 11600
rect 22277 11595 22343 11598
rect 23200 11568 24000 11598
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 0 11250 800 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 800 11190
rect 1577 11187 1643 11190
rect 23200 11024 24000 11144
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 0 10480 800 10600
rect 22277 10570 22343 10573
rect 23200 10570 24000 10600
rect 22277 10568 24000 10570
rect 22277 10512 22282 10568
rect 22338 10512 24000 10568
rect 22277 10510 24000 10512
rect 22277 10507 22343 10510
rect 23200 10480 24000 10510
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 22277 10026 22343 10029
rect 23200 10026 24000 10056
rect 22277 10024 24000 10026
rect 22277 9968 22282 10024
rect 22338 9968 24000 10024
rect 22277 9966 24000 9968
rect 22277 9963 22343 9966
rect 23200 9936 24000 9966
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 23200 9392 24000 9512
rect 3660 9280 3976 9281
rect 0 9210 800 9240
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 22277 8938 22343 8941
rect 23200 8938 24000 8968
rect 22277 8936 24000 8938
rect 22277 8880 22282 8936
rect 22338 8880 24000 8936
rect 22277 8878 24000 8880
rect 22277 8875 22343 8878
rect 23200 8848 24000 8878
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 0 8440 800 8560
rect 22277 8394 22343 8397
rect 23200 8394 24000 8424
rect 22277 8392 24000 8394
rect 22277 8336 22282 8392
rect 22338 8336 24000 8392
rect 22277 8334 24000 8336
rect 22277 8331 22343 8334
rect 23200 8304 24000 8334
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 23200 7760 24000 7880
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 22277 7306 22343 7309
rect 23200 7306 24000 7336
rect 22277 7304 24000 7306
rect 22277 7248 22282 7304
rect 22338 7248 24000 7304
rect 22277 7246 24000 7248
rect 22277 7243 22343 7246
rect 23200 7216 24000 7246
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 22277 6762 22343 6765
rect 23200 6762 24000 6792
rect 22277 6760 24000 6762
rect 22277 6704 22282 6760
rect 22338 6704 24000 6760
rect 22277 6702 24000 6704
rect 22277 6699 22343 6702
rect 23200 6672 24000 6702
rect 6374 6560 6690 6561
rect 0 6400 800 6520
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 23200 6128 24000 6248
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 22277 5674 22343 5677
rect 23200 5674 24000 5704
rect 22277 5672 24000 5674
rect 22277 5616 22282 5672
rect 22338 5616 24000 5672
rect 22277 5614 24000 5616
rect 22277 5611 22343 5614
rect 23200 5584 24000 5614
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 22277 5130 22343 5133
rect 23200 5130 24000 5160
rect 22277 5128 24000 5130
rect 22277 5072 22282 5128
rect 22338 5072 24000 5128
rect 22277 5070 24000 5072
rect 22277 5067 22343 5070
rect 23200 5040 24000 5070
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 23200 4496 24000 4616
rect 0 4360 800 4480
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 22277 4042 22343 4045
rect 23200 4042 24000 4072
rect 22277 4040 24000 4042
rect 22277 3984 22282 4040
rect 22338 3984 24000 4040
rect 22277 3982 24000 3984
rect 22277 3979 22343 3982
rect 23200 3952 24000 3982
rect 3660 3840 3976 3841
rect 0 3770 800 3800
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 22277 3498 22343 3501
rect 23200 3498 24000 3528
rect 22277 3496 24000 3498
rect 22277 3440 22282 3496
rect 22338 3440 24000 3496
rect 22277 3438 24000 3440
rect 22277 3435 22343 3438
rect 23200 3408 24000 3438
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 23200 2864 24000 2984
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 0 2320 800 2440
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
rect 0 1730 800 1760
rect 1577 1730 1643 1733
rect 0 1728 1643 1730
rect 0 1672 1582 1728
rect 1638 1672 1643 1728
rect 0 1670 1643 1672
rect 0 1640 800 1670
rect 1577 1667 1643 1670
rect 0 1050 800 1080
rect 1393 1050 1459 1053
rect 0 1048 1459 1050
rect 0 992 1398 1048
rect 1454 992 1459 1048
rect 0 990 1459 992
rect 0 960 800 990
rect 1393 987 1459 990
<< via3 >>
rect 3666 27772 3730 27776
rect 3666 27716 3670 27772
rect 3670 27716 3726 27772
rect 3726 27716 3730 27772
rect 3666 27712 3730 27716
rect 3746 27772 3810 27776
rect 3746 27716 3750 27772
rect 3750 27716 3806 27772
rect 3806 27716 3810 27772
rect 3746 27712 3810 27716
rect 3826 27772 3890 27776
rect 3826 27716 3830 27772
rect 3830 27716 3886 27772
rect 3886 27716 3890 27772
rect 3826 27712 3890 27716
rect 3906 27772 3970 27776
rect 3906 27716 3910 27772
rect 3910 27716 3966 27772
rect 3966 27716 3970 27772
rect 3906 27712 3970 27716
rect 9094 27772 9158 27776
rect 9094 27716 9098 27772
rect 9098 27716 9154 27772
rect 9154 27716 9158 27772
rect 9094 27712 9158 27716
rect 9174 27772 9238 27776
rect 9174 27716 9178 27772
rect 9178 27716 9234 27772
rect 9234 27716 9238 27772
rect 9174 27712 9238 27716
rect 9254 27772 9318 27776
rect 9254 27716 9258 27772
rect 9258 27716 9314 27772
rect 9314 27716 9318 27772
rect 9254 27712 9318 27716
rect 9334 27772 9398 27776
rect 9334 27716 9338 27772
rect 9338 27716 9394 27772
rect 9394 27716 9398 27772
rect 9334 27712 9398 27716
rect 14522 27772 14586 27776
rect 14522 27716 14526 27772
rect 14526 27716 14582 27772
rect 14582 27716 14586 27772
rect 14522 27712 14586 27716
rect 14602 27772 14666 27776
rect 14602 27716 14606 27772
rect 14606 27716 14662 27772
rect 14662 27716 14666 27772
rect 14602 27712 14666 27716
rect 14682 27772 14746 27776
rect 14682 27716 14686 27772
rect 14686 27716 14742 27772
rect 14742 27716 14746 27772
rect 14682 27712 14746 27716
rect 14762 27772 14826 27776
rect 14762 27716 14766 27772
rect 14766 27716 14822 27772
rect 14822 27716 14826 27772
rect 14762 27712 14826 27716
rect 19950 27772 20014 27776
rect 19950 27716 19954 27772
rect 19954 27716 20010 27772
rect 20010 27716 20014 27772
rect 19950 27712 20014 27716
rect 20030 27772 20094 27776
rect 20030 27716 20034 27772
rect 20034 27716 20090 27772
rect 20090 27716 20094 27772
rect 20030 27712 20094 27716
rect 20110 27772 20174 27776
rect 20110 27716 20114 27772
rect 20114 27716 20170 27772
rect 20170 27716 20174 27772
rect 20110 27712 20174 27716
rect 20190 27772 20254 27776
rect 20190 27716 20194 27772
rect 20194 27716 20250 27772
rect 20250 27716 20254 27772
rect 20190 27712 20254 27716
rect 6380 27228 6444 27232
rect 6380 27172 6384 27228
rect 6384 27172 6440 27228
rect 6440 27172 6444 27228
rect 6380 27168 6444 27172
rect 6460 27228 6524 27232
rect 6460 27172 6464 27228
rect 6464 27172 6520 27228
rect 6520 27172 6524 27228
rect 6460 27168 6524 27172
rect 6540 27228 6604 27232
rect 6540 27172 6544 27228
rect 6544 27172 6600 27228
rect 6600 27172 6604 27228
rect 6540 27168 6604 27172
rect 6620 27228 6684 27232
rect 6620 27172 6624 27228
rect 6624 27172 6680 27228
rect 6680 27172 6684 27228
rect 6620 27168 6684 27172
rect 11808 27228 11872 27232
rect 11808 27172 11812 27228
rect 11812 27172 11868 27228
rect 11868 27172 11872 27228
rect 11808 27168 11872 27172
rect 11888 27228 11952 27232
rect 11888 27172 11892 27228
rect 11892 27172 11948 27228
rect 11948 27172 11952 27228
rect 11888 27168 11952 27172
rect 11968 27228 12032 27232
rect 11968 27172 11972 27228
rect 11972 27172 12028 27228
rect 12028 27172 12032 27228
rect 11968 27168 12032 27172
rect 12048 27228 12112 27232
rect 12048 27172 12052 27228
rect 12052 27172 12108 27228
rect 12108 27172 12112 27228
rect 12048 27168 12112 27172
rect 17236 27228 17300 27232
rect 17236 27172 17240 27228
rect 17240 27172 17296 27228
rect 17296 27172 17300 27228
rect 17236 27168 17300 27172
rect 17316 27228 17380 27232
rect 17316 27172 17320 27228
rect 17320 27172 17376 27228
rect 17376 27172 17380 27228
rect 17316 27168 17380 27172
rect 17396 27228 17460 27232
rect 17396 27172 17400 27228
rect 17400 27172 17456 27228
rect 17456 27172 17460 27228
rect 17396 27168 17460 27172
rect 17476 27228 17540 27232
rect 17476 27172 17480 27228
rect 17480 27172 17536 27228
rect 17536 27172 17540 27228
rect 17476 27168 17540 27172
rect 22664 27228 22728 27232
rect 22664 27172 22668 27228
rect 22668 27172 22724 27228
rect 22724 27172 22728 27228
rect 22664 27168 22728 27172
rect 22744 27228 22808 27232
rect 22744 27172 22748 27228
rect 22748 27172 22804 27228
rect 22804 27172 22808 27228
rect 22744 27168 22808 27172
rect 22824 27228 22888 27232
rect 22824 27172 22828 27228
rect 22828 27172 22884 27228
rect 22884 27172 22888 27228
rect 22824 27168 22888 27172
rect 22904 27228 22968 27232
rect 22904 27172 22908 27228
rect 22908 27172 22964 27228
rect 22964 27172 22968 27228
rect 22904 27168 22968 27172
rect 3666 26684 3730 26688
rect 3666 26628 3670 26684
rect 3670 26628 3726 26684
rect 3726 26628 3730 26684
rect 3666 26624 3730 26628
rect 3746 26684 3810 26688
rect 3746 26628 3750 26684
rect 3750 26628 3806 26684
rect 3806 26628 3810 26684
rect 3746 26624 3810 26628
rect 3826 26684 3890 26688
rect 3826 26628 3830 26684
rect 3830 26628 3886 26684
rect 3886 26628 3890 26684
rect 3826 26624 3890 26628
rect 3906 26684 3970 26688
rect 3906 26628 3910 26684
rect 3910 26628 3966 26684
rect 3966 26628 3970 26684
rect 3906 26624 3970 26628
rect 9094 26684 9158 26688
rect 9094 26628 9098 26684
rect 9098 26628 9154 26684
rect 9154 26628 9158 26684
rect 9094 26624 9158 26628
rect 9174 26684 9238 26688
rect 9174 26628 9178 26684
rect 9178 26628 9234 26684
rect 9234 26628 9238 26684
rect 9174 26624 9238 26628
rect 9254 26684 9318 26688
rect 9254 26628 9258 26684
rect 9258 26628 9314 26684
rect 9314 26628 9318 26684
rect 9254 26624 9318 26628
rect 9334 26684 9398 26688
rect 9334 26628 9338 26684
rect 9338 26628 9394 26684
rect 9394 26628 9398 26684
rect 9334 26624 9398 26628
rect 14522 26684 14586 26688
rect 14522 26628 14526 26684
rect 14526 26628 14582 26684
rect 14582 26628 14586 26684
rect 14522 26624 14586 26628
rect 14602 26684 14666 26688
rect 14602 26628 14606 26684
rect 14606 26628 14662 26684
rect 14662 26628 14666 26684
rect 14602 26624 14666 26628
rect 14682 26684 14746 26688
rect 14682 26628 14686 26684
rect 14686 26628 14742 26684
rect 14742 26628 14746 26684
rect 14682 26624 14746 26628
rect 14762 26684 14826 26688
rect 14762 26628 14766 26684
rect 14766 26628 14822 26684
rect 14822 26628 14826 26684
rect 14762 26624 14826 26628
rect 19950 26684 20014 26688
rect 19950 26628 19954 26684
rect 19954 26628 20010 26684
rect 20010 26628 20014 26684
rect 19950 26624 20014 26628
rect 20030 26684 20094 26688
rect 20030 26628 20034 26684
rect 20034 26628 20090 26684
rect 20090 26628 20094 26684
rect 20030 26624 20094 26628
rect 20110 26684 20174 26688
rect 20110 26628 20114 26684
rect 20114 26628 20170 26684
rect 20170 26628 20174 26684
rect 20110 26624 20174 26628
rect 20190 26684 20254 26688
rect 20190 26628 20194 26684
rect 20194 26628 20250 26684
rect 20250 26628 20254 26684
rect 20190 26624 20254 26628
rect 6380 26140 6444 26144
rect 6380 26084 6384 26140
rect 6384 26084 6440 26140
rect 6440 26084 6444 26140
rect 6380 26080 6444 26084
rect 6460 26140 6524 26144
rect 6460 26084 6464 26140
rect 6464 26084 6520 26140
rect 6520 26084 6524 26140
rect 6460 26080 6524 26084
rect 6540 26140 6604 26144
rect 6540 26084 6544 26140
rect 6544 26084 6600 26140
rect 6600 26084 6604 26140
rect 6540 26080 6604 26084
rect 6620 26140 6684 26144
rect 6620 26084 6624 26140
rect 6624 26084 6680 26140
rect 6680 26084 6684 26140
rect 6620 26080 6684 26084
rect 11808 26140 11872 26144
rect 11808 26084 11812 26140
rect 11812 26084 11868 26140
rect 11868 26084 11872 26140
rect 11808 26080 11872 26084
rect 11888 26140 11952 26144
rect 11888 26084 11892 26140
rect 11892 26084 11948 26140
rect 11948 26084 11952 26140
rect 11888 26080 11952 26084
rect 11968 26140 12032 26144
rect 11968 26084 11972 26140
rect 11972 26084 12028 26140
rect 12028 26084 12032 26140
rect 11968 26080 12032 26084
rect 12048 26140 12112 26144
rect 12048 26084 12052 26140
rect 12052 26084 12108 26140
rect 12108 26084 12112 26140
rect 12048 26080 12112 26084
rect 17236 26140 17300 26144
rect 17236 26084 17240 26140
rect 17240 26084 17296 26140
rect 17296 26084 17300 26140
rect 17236 26080 17300 26084
rect 17316 26140 17380 26144
rect 17316 26084 17320 26140
rect 17320 26084 17376 26140
rect 17376 26084 17380 26140
rect 17316 26080 17380 26084
rect 17396 26140 17460 26144
rect 17396 26084 17400 26140
rect 17400 26084 17456 26140
rect 17456 26084 17460 26140
rect 17396 26080 17460 26084
rect 17476 26140 17540 26144
rect 17476 26084 17480 26140
rect 17480 26084 17536 26140
rect 17536 26084 17540 26140
rect 17476 26080 17540 26084
rect 22664 26140 22728 26144
rect 22664 26084 22668 26140
rect 22668 26084 22724 26140
rect 22724 26084 22728 26140
rect 22664 26080 22728 26084
rect 22744 26140 22808 26144
rect 22744 26084 22748 26140
rect 22748 26084 22804 26140
rect 22804 26084 22808 26140
rect 22744 26080 22808 26084
rect 22824 26140 22888 26144
rect 22824 26084 22828 26140
rect 22828 26084 22884 26140
rect 22884 26084 22888 26140
rect 22824 26080 22888 26084
rect 22904 26140 22968 26144
rect 22904 26084 22908 26140
rect 22908 26084 22964 26140
rect 22964 26084 22968 26140
rect 22904 26080 22968 26084
rect 3666 25596 3730 25600
rect 3666 25540 3670 25596
rect 3670 25540 3726 25596
rect 3726 25540 3730 25596
rect 3666 25536 3730 25540
rect 3746 25596 3810 25600
rect 3746 25540 3750 25596
rect 3750 25540 3806 25596
rect 3806 25540 3810 25596
rect 3746 25536 3810 25540
rect 3826 25596 3890 25600
rect 3826 25540 3830 25596
rect 3830 25540 3886 25596
rect 3886 25540 3890 25596
rect 3826 25536 3890 25540
rect 3906 25596 3970 25600
rect 3906 25540 3910 25596
rect 3910 25540 3966 25596
rect 3966 25540 3970 25596
rect 3906 25536 3970 25540
rect 9094 25596 9158 25600
rect 9094 25540 9098 25596
rect 9098 25540 9154 25596
rect 9154 25540 9158 25596
rect 9094 25536 9158 25540
rect 9174 25596 9238 25600
rect 9174 25540 9178 25596
rect 9178 25540 9234 25596
rect 9234 25540 9238 25596
rect 9174 25536 9238 25540
rect 9254 25596 9318 25600
rect 9254 25540 9258 25596
rect 9258 25540 9314 25596
rect 9314 25540 9318 25596
rect 9254 25536 9318 25540
rect 9334 25596 9398 25600
rect 9334 25540 9338 25596
rect 9338 25540 9394 25596
rect 9394 25540 9398 25596
rect 9334 25536 9398 25540
rect 14522 25596 14586 25600
rect 14522 25540 14526 25596
rect 14526 25540 14582 25596
rect 14582 25540 14586 25596
rect 14522 25536 14586 25540
rect 14602 25596 14666 25600
rect 14602 25540 14606 25596
rect 14606 25540 14662 25596
rect 14662 25540 14666 25596
rect 14602 25536 14666 25540
rect 14682 25596 14746 25600
rect 14682 25540 14686 25596
rect 14686 25540 14742 25596
rect 14742 25540 14746 25596
rect 14682 25536 14746 25540
rect 14762 25596 14826 25600
rect 14762 25540 14766 25596
rect 14766 25540 14822 25596
rect 14822 25540 14826 25596
rect 14762 25536 14826 25540
rect 19950 25596 20014 25600
rect 19950 25540 19954 25596
rect 19954 25540 20010 25596
rect 20010 25540 20014 25596
rect 19950 25536 20014 25540
rect 20030 25596 20094 25600
rect 20030 25540 20034 25596
rect 20034 25540 20090 25596
rect 20090 25540 20094 25596
rect 20030 25536 20094 25540
rect 20110 25596 20174 25600
rect 20110 25540 20114 25596
rect 20114 25540 20170 25596
rect 20170 25540 20174 25596
rect 20110 25536 20174 25540
rect 20190 25596 20254 25600
rect 20190 25540 20194 25596
rect 20194 25540 20250 25596
rect 20250 25540 20254 25596
rect 20190 25536 20254 25540
rect 6380 25052 6444 25056
rect 6380 24996 6384 25052
rect 6384 24996 6440 25052
rect 6440 24996 6444 25052
rect 6380 24992 6444 24996
rect 6460 25052 6524 25056
rect 6460 24996 6464 25052
rect 6464 24996 6520 25052
rect 6520 24996 6524 25052
rect 6460 24992 6524 24996
rect 6540 25052 6604 25056
rect 6540 24996 6544 25052
rect 6544 24996 6600 25052
rect 6600 24996 6604 25052
rect 6540 24992 6604 24996
rect 6620 25052 6684 25056
rect 6620 24996 6624 25052
rect 6624 24996 6680 25052
rect 6680 24996 6684 25052
rect 6620 24992 6684 24996
rect 11808 25052 11872 25056
rect 11808 24996 11812 25052
rect 11812 24996 11868 25052
rect 11868 24996 11872 25052
rect 11808 24992 11872 24996
rect 11888 25052 11952 25056
rect 11888 24996 11892 25052
rect 11892 24996 11948 25052
rect 11948 24996 11952 25052
rect 11888 24992 11952 24996
rect 11968 25052 12032 25056
rect 11968 24996 11972 25052
rect 11972 24996 12028 25052
rect 12028 24996 12032 25052
rect 11968 24992 12032 24996
rect 12048 25052 12112 25056
rect 12048 24996 12052 25052
rect 12052 24996 12108 25052
rect 12108 24996 12112 25052
rect 12048 24992 12112 24996
rect 17236 25052 17300 25056
rect 17236 24996 17240 25052
rect 17240 24996 17296 25052
rect 17296 24996 17300 25052
rect 17236 24992 17300 24996
rect 17316 25052 17380 25056
rect 17316 24996 17320 25052
rect 17320 24996 17376 25052
rect 17376 24996 17380 25052
rect 17316 24992 17380 24996
rect 17396 25052 17460 25056
rect 17396 24996 17400 25052
rect 17400 24996 17456 25052
rect 17456 24996 17460 25052
rect 17396 24992 17460 24996
rect 17476 25052 17540 25056
rect 17476 24996 17480 25052
rect 17480 24996 17536 25052
rect 17536 24996 17540 25052
rect 17476 24992 17540 24996
rect 22664 25052 22728 25056
rect 22664 24996 22668 25052
rect 22668 24996 22724 25052
rect 22724 24996 22728 25052
rect 22664 24992 22728 24996
rect 22744 25052 22808 25056
rect 22744 24996 22748 25052
rect 22748 24996 22804 25052
rect 22804 24996 22808 25052
rect 22744 24992 22808 24996
rect 22824 25052 22888 25056
rect 22824 24996 22828 25052
rect 22828 24996 22884 25052
rect 22884 24996 22888 25052
rect 22824 24992 22888 24996
rect 22904 25052 22968 25056
rect 22904 24996 22908 25052
rect 22908 24996 22964 25052
rect 22964 24996 22968 25052
rect 22904 24992 22968 24996
rect 3666 24508 3730 24512
rect 3666 24452 3670 24508
rect 3670 24452 3726 24508
rect 3726 24452 3730 24508
rect 3666 24448 3730 24452
rect 3746 24508 3810 24512
rect 3746 24452 3750 24508
rect 3750 24452 3806 24508
rect 3806 24452 3810 24508
rect 3746 24448 3810 24452
rect 3826 24508 3890 24512
rect 3826 24452 3830 24508
rect 3830 24452 3886 24508
rect 3886 24452 3890 24508
rect 3826 24448 3890 24452
rect 3906 24508 3970 24512
rect 3906 24452 3910 24508
rect 3910 24452 3966 24508
rect 3966 24452 3970 24508
rect 3906 24448 3970 24452
rect 9094 24508 9158 24512
rect 9094 24452 9098 24508
rect 9098 24452 9154 24508
rect 9154 24452 9158 24508
rect 9094 24448 9158 24452
rect 9174 24508 9238 24512
rect 9174 24452 9178 24508
rect 9178 24452 9234 24508
rect 9234 24452 9238 24508
rect 9174 24448 9238 24452
rect 9254 24508 9318 24512
rect 9254 24452 9258 24508
rect 9258 24452 9314 24508
rect 9314 24452 9318 24508
rect 9254 24448 9318 24452
rect 9334 24508 9398 24512
rect 9334 24452 9338 24508
rect 9338 24452 9394 24508
rect 9394 24452 9398 24508
rect 9334 24448 9398 24452
rect 14522 24508 14586 24512
rect 14522 24452 14526 24508
rect 14526 24452 14582 24508
rect 14582 24452 14586 24508
rect 14522 24448 14586 24452
rect 14602 24508 14666 24512
rect 14602 24452 14606 24508
rect 14606 24452 14662 24508
rect 14662 24452 14666 24508
rect 14602 24448 14666 24452
rect 14682 24508 14746 24512
rect 14682 24452 14686 24508
rect 14686 24452 14742 24508
rect 14742 24452 14746 24508
rect 14682 24448 14746 24452
rect 14762 24508 14826 24512
rect 14762 24452 14766 24508
rect 14766 24452 14822 24508
rect 14822 24452 14826 24508
rect 14762 24448 14826 24452
rect 19950 24508 20014 24512
rect 19950 24452 19954 24508
rect 19954 24452 20010 24508
rect 20010 24452 20014 24508
rect 19950 24448 20014 24452
rect 20030 24508 20094 24512
rect 20030 24452 20034 24508
rect 20034 24452 20090 24508
rect 20090 24452 20094 24508
rect 20030 24448 20094 24452
rect 20110 24508 20174 24512
rect 20110 24452 20114 24508
rect 20114 24452 20170 24508
rect 20170 24452 20174 24508
rect 20110 24448 20174 24452
rect 20190 24508 20254 24512
rect 20190 24452 20194 24508
rect 20194 24452 20250 24508
rect 20250 24452 20254 24508
rect 20190 24448 20254 24452
rect 6380 23964 6444 23968
rect 6380 23908 6384 23964
rect 6384 23908 6440 23964
rect 6440 23908 6444 23964
rect 6380 23904 6444 23908
rect 6460 23964 6524 23968
rect 6460 23908 6464 23964
rect 6464 23908 6520 23964
rect 6520 23908 6524 23964
rect 6460 23904 6524 23908
rect 6540 23964 6604 23968
rect 6540 23908 6544 23964
rect 6544 23908 6600 23964
rect 6600 23908 6604 23964
rect 6540 23904 6604 23908
rect 6620 23964 6684 23968
rect 6620 23908 6624 23964
rect 6624 23908 6680 23964
rect 6680 23908 6684 23964
rect 6620 23904 6684 23908
rect 11808 23964 11872 23968
rect 11808 23908 11812 23964
rect 11812 23908 11868 23964
rect 11868 23908 11872 23964
rect 11808 23904 11872 23908
rect 11888 23964 11952 23968
rect 11888 23908 11892 23964
rect 11892 23908 11948 23964
rect 11948 23908 11952 23964
rect 11888 23904 11952 23908
rect 11968 23964 12032 23968
rect 11968 23908 11972 23964
rect 11972 23908 12028 23964
rect 12028 23908 12032 23964
rect 11968 23904 12032 23908
rect 12048 23964 12112 23968
rect 12048 23908 12052 23964
rect 12052 23908 12108 23964
rect 12108 23908 12112 23964
rect 12048 23904 12112 23908
rect 17236 23964 17300 23968
rect 17236 23908 17240 23964
rect 17240 23908 17296 23964
rect 17296 23908 17300 23964
rect 17236 23904 17300 23908
rect 17316 23964 17380 23968
rect 17316 23908 17320 23964
rect 17320 23908 17376 23964
rect 17376 23908 17380 23964
rect 17316 23904 17380 23908
rect 17396 23964 17460 23968
rect 17396 23908 17400 23964
rect 17400 23908 17456 23964
rect 17456 23908 17460 23964
rect 17396 23904 17460 23908
rect 17476 23964 17540 23968
rect 17476 23908 17480 23964
rect 17480 23908 17536 23964
rect 17536 23908 17540 23964
rect 17476 23904 17540 23908
rect 22664 23964 22728 23968
rect 22664 23908 22668 23964
rect 22668 23908 22724 23964
rect 22724 23908 22728 23964
rect 22664 23904 22728 23908
rect 22744 23964 22808 23968
rect 22744 23908 22748 23964
rect 22748 23908 22804 23964
rect 22804 23908 22808 23964
rect 22744 23904 22808 23908
rect 22824 23964 22888 23968
rect 22824 23908 22828 23964
rect 22828 23908 22884 23964
rect 22884 23908 22888 23964
rect 22824 23904 22888 23908
rect 22904 23964 22968 23968
rect 22904 23908 22908 23964
rect 22908 23908 22964 23964
rect 22964 23908 22968 23964
rect 22904 23904 22968 23908
rect 3666 23420 3730 23424
rect 3666 23364 3670 23420
rect 3670 23364 3726 23420
rect 3726 23364 3730 23420
rect 3666 23360 3730 23364
rect 3746 23420 3810 23424
rect 3746 23364 3750 23420
rect 3750 23364 3806 23420
rect 3806 23364 3810 23420
rect 3746 23360 3810 23364
rect 3826 23420 3890 23424
rect 3826 23364 3830 23420
rect 3830 23364 3886 23420
rect 3886 23364 3890 23420
rect 3826 23360 3890 23364
rect 3906 23420 3970 23424
rect 3906 23364 3910 23420
rect 3910 23364 3966 23420
rect 3966 23364 3970 23420
rect 3906 23360 3970 23364
rect 9094 23420 9158 23424
rect 9094 23364 9098 23420
rect 9098 23364 9154 23420
rect 9154 23364 9158 23420
rect 9094 23360 9158 23364
rect 9174 23420 9238 23424
rect 9174 23364 9178 23420
rect 9178 23364 9234 23420
rect 9234 23364 9238 23420
rect 9174 23360 9238 23364
rect 9254 23420 9318 23424
rect 9254 23364 9258 23420
rect 9258 23364 9314 23420
rect 9314 23364 9318 23420
rect 9254 23360 9318 23364
rect 9334 23420 9398 23424
rect 9334 23364 9338 23420
rect 9338 23364 9394 23420
rect 9394 23364 9398 23420
rect 9334 23360 9398 23364
rect 14522 23420 14586 23424
rect 14522 23364 14526 23420
rect 14526 23364 14582 23420
rect 14582 23364 14586 23420
rect 14522 23360 14586 23364
rect 14602 23420 14666 23424
rect 14602 23364 14606 23420
rect 14606 23364 14662 23420
rect 14662 23364 14666 23420
rect 14602 23360 14666 23364
rect 14682 23420 14746 23424
rect 14682 23364 14686 23420
rect 14686 23364 14742 23420
rect 14742 23364 14746 23420
rect 14682 23360 14746 23364
rect 14762 23420 14826 23424
rect 14762 23364 14766 23420
rect 14766 23364 14822 23420
rect 14822 23364 14826 23420
rect 14762 23360 14826 23364
rect 19950 23420 20014 23424
rect 19950 23364 19954 23420
rect 19954 23364 20010 23420
rect 20010 23364 20014 23420
rect 19950 23360 20014 23364
rect 20030 23420 20094 23424
rect 20030 23364 20034 23420
rect 20034 23364 20090 23420
rect 20090 23364 20094 23420
rect 20030 23360 20094 23364
rect 20110 23420 20174 23424
rect 20110 23364 20114 23420
rect 20114 23364 20170 23420
rect 20170 23364 20174 23420
rect 20110 23360 20174 23364
rect 20190 23420 20254 23424
rect 20190 23364 20194 23420
rect 20194 23364 20250 23420
rect 20250 23364 20254 23420
rect 20190 23360 20254 23364
rect 6380 22876 6444 22880
rect 6380 22820 6384 22876
rect 6384 22820 6440 22876
rect 6440 22820 6444 22876
rect 6380 22816 6444 22820
rect 6460 22876 6524 22880
rect 6460 22820 6464 22876
rect 6464 22820 6520 22876
rect 6520 22820 6524 22876
rect 6460 22816 6524 22820
rect 6540 22876 6604 22880
rect 6540 22820 6544 22876
rect 6544 22820 6600 22876
rect 6600 22820 6604 22876
rect 6540 22816 6604 22820
rect 6620 22876 6684 22880
rect 6620 22820 6624 22876
rect 6624 22820 6680 22876
rect 6680 22820 6684 22876
rect 6620 22816 6684 22820
rect 11808 22876 11872 22880
rect 11808 22820 11812 22876
rect 11812 22820 11868 22876
rect 11868 22820 11872 22876
rect 11808 22816 11872 22820
rect 11888 22876 11952 22880
rect 11888 22820 11892 22876
rect 11892 22820 11948 22876
rect 11948 22820 11952 22876
rect 11888 22816 11952 22820
rect 11968 22876 12032 22880
rect 11968 22820 11972 22876
rect 11972 22820 12028 22876
rect 12028 22820 12032 22876
rect 11968 22816 12032 22820
rect 12048 22876 12112 22880
rect 12048 22820 12052 22876
rect 12052 22820 12108 22876
rect 12108 22820 12112 22876
rect 12048 22816 12112 22820
rect 17236 22876 17300 22880
rect 17236 22820 17240 22876
rect 17240 22820 17296 22876
rect 17296 22820 17300 22876
rect 17236 22816 17300 22820
rect 17316 22876 17380 22880
rect 17316 22820 17320 22876
rect 17320 22820 17376 22876
rect 17376 22820 17380 22876
rect 17316 22816 17380 22820
rect 17396 22876 17460 22880
rect 17396 22820 17400 22876
rect 17400 22820 17456 22876
rect 17456 22820 17460 22876
rect 17396 22816 17460 22820
rect 17476 22876 17540 22880
rect 17476 22820 17480 22876
rect 17480 22820 17536 22876
rect 17536 22820 17540 22876
rect 17476 22816 17540 22820
rect 22664 22876 22728 22880
rect 22664 22820 22668 22876
rect 22668 22820 22724 22876
rect 22724 22820 22728 22876
rect 22664 22816 22728 22820
rect 22744 22876 22808 22880
rect 22744 22820 22748 22876
rect 22748 22820 22804 22876
rect 22804 22820 22808 22876
rect 22744 22816 22808 22820
rect 22824 22876 22888 22880
rect 22824 22820 22828 22876
rect 22828 22820 22884 22876
rect 22884 22820 22888 22876
rect 22824 22816 22888 22820
rect 22904 22876 22968 22880
rect 22904 22820 22908 22876
rect 22908 22820 22964 22876
rect 22964 22820 22968 22876
rect 22904 22816 22968 22820
rect 3666 22332 3730 22336
rect 3666 22276 3670 22332
rect 3670 22276 3726 22332
rect 3726 22276 3730 22332
rect 3666 22272 3730 22276
rect 3746 22332 3810 22336
rect 3746 22276 3750 22332
rect 3750 22276 3806 22332
rect 3806 22276 3810 22332
rect 3746 22272 3810 22276
rect 3826 22332 3890 22336
rect 3826 22276 3830 22332
rect 3830 22276 3886 22332
rect 3886 22276 3890 22332
rect 3826 22272 3890 22276
rect 3906 22332 3970 22336
rect 3906 22276 3910 22332
rect 3910 22276 3966 22332
rect 3966 22276 3970 22332
rect 3906 22272 3970 22276
rect 9094 22332 9158 22336
rect 9094 22276 9098 22332
rect 9098 22276 9154 22332
rect 9154 22276 9158 22332
rect 9094 22272 9158 22276
rect 9174 22332 9238 22336
rect 9174 22276 9178 22332
rect 9178 22276 9234 22332
rect 9234 22276 9238 22332
rect 9174 22272 9238 22276
rect 9254 22332 9318 22336
rect 9254 22276 9258 22332
rect 9258 22276 9314 22332
rect 9314 22276 9318 22332
rect 9254 22272 9318 22276
rect 9334 22332 9398 22336
rect 9334 22276 9338 22332
rect 9338 22276 9394 22332
rect 9394 22276 9398 22332
rect 9334 22272 9398 22276
rect 14522 22332 14586 22336
rect 14522 22276 14526 22332
rect 14526 22276 14582 22332
rect 14582 22276 14586 22332
rect 14522 22272 14586 22276
rect 14602 22332 14666 22336
rect 14602 22276 14606 22332
rect 14606 22276 14662 22332
rect 14662 22276 14666 22332
rect 14602 22272 14666 22276
rect 14682 22332 14746 22336
rect 14682 22276 14686 22332
rect 14686 22276 14742 22332
rect 14742 22276 14746 22332
rect 14682 22272 14746 22276
rect 14762 22332 14826 22336
rect 14762 22276 14766 22332
rect 14766 22276 14822 22332
rect 14822 22276 14826 22332
rect 14762 22272 14826 22276
rect 19950 22332 20014 22336
rect 19950 22276 19954 22332
rect 19954 22276 20010 22332
rect 20010 22276 20014 22332
rect 19950 22272 20014 22276
rect 20030 22332 20094 22336
rect 20030 22276 20034 22332
rect 20034 22276 20090 22332
rect 20090 22276 20094 22332
rect 20030 22272 20094 22276
rect 20110 22332 20174 22336
rect 20110 22276 20114 22332
rect 20114 22276 20170 22332
rect 20170 22276 20174 22332
rect 20110 22272 20174 22276
rect 20190 22332 20254 22336
rect 20190 22276 20194 22332
rect 20194 22276 20250 22332
rect 20250 22276 20254 22332
rect 20190 22272 20254 22276
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 27776 3978 27792
rect 3658 27712 3666 27776
rect 3730 27712 3746 27776
rect 3810 27712 3826 27776
rect 3890 27712 3906 27776
rect 3970 27712 3978 27776
rect 3658 26688 3978 27712
rect 3658 26624 3666 26688
rect 3730 26624 3746 26688
rect 3810 26624 3826 26688
rect 3890 26624 3906 26688
rect 3970 26624 3978 26688
rect 3658 25600 3978 26624
rect 3658 25536 3666 25600
rect 3730 25536 3746 25600
rect 3810 25536 3826 25600
rect 3890 25536 3906 25600
rect 3970 25536 3978 25600
rect 3658 24512 3978 25536
rect 3658 24448 3666 24512
rect 3730 24448 3746 24512
rect 3810 24448 3826 24512
rect 3890 24448 3906 24512
rect 3970 24448 3978 24512
rect 3658 23424 3978 24448
rect 3658 23360 3666 23424
rect 3730 23360 3746 23424
rect 3810 23360 3826 23424
rect 3890 23360 3906 23424
rect 3970 23360 3978 23424
rect 3658 22336 3978 23360
rect 3658 22272 3666 22336
rect 3730 22272 3746 22336
rect 3810 22272 3826 22336
rect 3890 22272 3906 22336
rect 3970 22272 3978 22336
rect 3658 21248 3978 22272
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 27232 6692 27792
rect 6372 27168 6380 27232
rect 6444 27168 6460 27232
rect 6524 27168 6540 27232
rect 6604 27168 6620 27232
rect 6684 27168 6692 27232
rect 6372 26144 6692 27168
rect 6372 26080 6380 26144
rect 6444 26080 6460 26144
rect 6524 26080 6540 26144
rect 6604 26080 6620 26144
rect 6684 26080 6692 26144
rect 6372 25056 6692 26080
rect 6372 24992 6380 25056
rect 6444 24992 6460 25056
rect 6524 24992 6540 25056
rect 6604 24992 6620 25056
rect 6684 24992 6692 25056
rect 6372 23968 6692 24992
rect 6372 23904 6380 23968
rect 6444 23904 6460 23968
rect 6524 23904 6540 23968
rect 6604 23904 6620 23968
rect 6684 23904 6692 23968
rect 6372 22880 6692 23904
rect 6372 22816 6380 22880
rect 6444 22816 6460 22880
rect 6524 22816 6540 22880
rect 6604 22816 6620 22880
rect 6684 22816 6692 22880
rect 6372 21792 6692 22816
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 27776 9406 27792
rect 9086 27712 9094 27776
rect 9158 27712 9174 27776
rect 9238 27712 9254 27776
rect 9318 27712 9334 27776
rect 9398 27712 9406 27776
rect 9086 26688 9406 27712
rect 9086 26624 9094 26688
rect 9158 26624 9174 26688
rect 9238 26624 9254 26688
rect 9318 26624 9334 26688
rect 9398 26624 9406 26688
rect 9086 25600 9406 26624
rect 9086 25536 9094 25600
rect 9158 25536 9174 25600
rect 9238 25536 9254 25600
rect 9318 25536 9334 25600
rect 9398 25536 9406 25600
rect 9086 24512 9406 25536
rect 9086 24448 9094 24512
rect 9158 24448 9174 24512
rect 9238 24448 9254 24512
rect 9318 24448 9334 24512
rect 9398 24448 9406 24512
rect 9086 23424 9406 24448
rect 9086 23360 9094 23424
rect 9158 23360 9174 23424
rect 9238 23360 9254 23424
rect 9318 23360 9334 23424
rect 9398 23360 9406 23424
rect 9086 22336 9406 23360
rect 9086 22272 9094 22336
rect 9158 22272 9174 22336
rect 9238 22272 9254 22336
rect 9318 22272 9334 22336
rect 9398 22272 9406 22336
rect 9086 21248 9406 22272
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 27232 12120 27792
rect 11800 27168 11808 27232
rect 11872 27168 11888 27232
rect 11952 27168 11968 27232
rect 12032 27168 12048 27232
rect 12112 27168 12120 27232
rect 11800 26144 12120 27168
rect 11800 26080 11808 26144
rect 11872 26080 11888 26144
rect 11952 26080 11968 26144
rect 12032 26080 12048 26144
rect 12112 26080 12120 26144
rect 11800 25056 12120 26080
rect 11800 24992 11808 25056
rect 11872 24992 11888 25056
rect 11952 24992 11968 25056
rect 12032 24992 12048 25056
rect 12112 24992 12120 25056
rect 11800 23968 12120 24992
rect 11800 23904 11808 23968
rect 11872 23904 11888 23968
rect 11952 23904 11968 23968
rect 12032 23904 12048 23968
rect 12112 23904 12120 23968
rect 11800 22880 12120 23904
rect 11800 22816 11808 22880
rect 11872 22816 11888 22880
rect 11952 22816 11968 22880
rect 12032 22816 12048 22880
rect 12112 22816 12120 22880
rect 11800 21792 12120 22816
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 27776 14834 27792
rect 14514 27712 14522 27776
rect 14586 27712 14602 27776
rect 14666 27712 14682 27776
rect 14746 27712 14762 27776
rect 14826 27712 14834 27776
rect 14514 26688 14834 27712
rect 14514 26624 14522 26688
rect 14586 26624 14602 26688
rect 14666 26624 14682 26688
rect 14746 26624 14762 26688
rect 14826 26624 14834 26688
rect 14514 25600 14834 26624
rect 14514 25536 14522 25600
rect 14586 25536 14602 25600
rect 14666 25536 14682 25600
rect 14746 25536 14762 25600
rect 14826 25536 14834 25600
rect 14514 24512 14834 25536
rect 14514 24448 14522 24512
rect 14586 24448 14602 24512
rect 14666 24448 14682 24512
rect 14746 24448 14762 24512
rect 14826 24448 14834 24512
rect 14514 23424 14834 24448
rect 14514 23360 14522 23424
rect 14586 23360 14602 23424
rect 14666 23360 14682 23424
rect 14746 23360 14762 23424
rect 14826 23360 14834 23424
rect 14514 22336 14834 23360
rect 14514 22272 14522 22336
rect 14586 22272 14602 22336
rect 14666 22272 14682 22336
rect 14746 22272 14762 22336
rect 14826 22272 14834 22336
rect 14514 21248 14834 22272
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 27232 17548 27792
rect 17228 27168 17236 27232
rect 17300 27168 17316 27232
rect 17380 27168 17396 27232
rect 17460 27168 17476 27232
rect 17540 27168 17548 27232
rect 17228 26144 17548 27168
rect 17228 26080 17236 26144
rect 17300 26080 17316 26144
rect 17380 26080 17396 26144
rect 17460 26080 17476 26144
rect 17540 26080 17548 26144
rect 17228 25056 17548 26080
rect 17228 24992 17236 25056
rect 17300 24992 17316 25056
rect 17380 24992 17396 25056
rect 17460 24992 17476 25056
rect 17540 24992 17548 25056
rect 17228 23968 17548 24992
rect 17228 23904 17236 23968
rect 17300 23904 17316 23968
rect 17380 23904 17396 23968
rect 17460 23904 17476 23968
rect 17540 23904 17548 23968
rect 17228 22880 17548 23904
rect 17228 22816 17236 22880
rect 17300 22816 17316 22880
rect 17380 22816 17396 22880
rect 17460 22816 17476 22880
rect 17540 22816 17548 22880
rect 17228 21792 17548 22816
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 27776 20262 27792
rect 19942 27712 19950 27776
rect 20014 27712 20030 27776
rect 20094 27712 20110 27776
rect 20174 27712 20190 27776
rect 20254 27712 20262 27776
rect 19942 26688 20262 27712
rect 19942 26624 19950 26688
rect 20014 26624 20030 26688
rect 20094 26624 20110 26688
rect 20174 26624 20190 26688
rect 20254 26624 20262 26688
rect 19942 25600 20262 26624
rect 19942 25536 19950 25600
rect 20014 25536 20030 25600
rect 20094 25536 20110 25600
rect 20174 25536 20190 25600
rect 20254 25536 20262 25600
rect 19942 24512 20262 25536
rect 19942 24448 19950 24512
rect 20014 24448 20030 24512
rect 20094 24448 20110 24512
rect 20174 24448 20190 24512
rect 20254 24448 20262 24512
rect 19942 23424 20262 24448
rect 19942 23360 19950 23424
rect 20014 23360 20030 23424
rect 20094 23360 20110 23424
rect 20174 23360 20190 23424
rect 20254 23360 20262 23424
rect 19942 22336 20262 23360
rect 19942 22272 19950 22336
rect 20014 22272 20030 22336
rect 20094 22272 20110 22336
rect 20174 22272 20190 22336
rect 20254 22272 20262 22336
rect 19942 21248 20262 22272
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 27232 22976 27792
rect 22656 27168 22664 27232
rect 22728 27168 22744 27232
rect 22808 27168 22824 27232
rect 22888 27168 22904 27232
rect 22968 27168 22976 27232
rect 22656 26144 22976 27168
rect 22656 26080 22664 26144
rect 22728 26080 22744 26144
rect 22808 26080 22824 26144
rect 22888 26080 22904 26144
rect 22968 26080 22976 26144
rect 22656 25056 22976 26080
rect 22656 24992 22664 25056
rect 22728 24992 22744 25056
rect 22808 24992 22824 25056
rect 22888 24992 22904 25056
rect 22968 24992 22976 25056
rect 22656 23968 22976 24992
rect 22656 23904 22664 23968
rect 22728 23904 22744 23968
rect 22808 23904 22824 23968
rect 22888 23904 22904 23968
rect 22968 23904 22976 23968
rect 22656 22880 22976 23904
rect 22656 22816 22664 22880
rect 22728 22816 22744 22880
rect 22808 22816 22824 22880
rect 22888 22816 22904 22880
rect 22968 22816 22976 22880
rect 22656 21792 22976 22816
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1666464484
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1666464484
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_231
timestamp 1666464484
transform 1 0 22356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1666464484
transform 1 0 22356 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_227
timestamp 1666464484
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_231
timestamp 1666464484
transform 1 0 22356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1666464484
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1666464484
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1666464484
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1666464484
transform 1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_231
timestamp 1666464484
transform 1 0 22356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 1666464484
transform 1 0 22356 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_231
timestamp 1666464484
transform 1 0 22356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_227
timestamp 1666464484
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1666464484
transform 1 0 22356 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 1666464484
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1666464484
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_227
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1666464484
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1666464484
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_231
timestamp 1666464484
transform 1 0 22356 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_231
timestamp 1666464484
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1666464484
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1666464484
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_231
timestamp 1666464484
transform 1 0 22356 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_227
timestamp 1666464484
transform 1 0 21988 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_231
timestamp 1666464484
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1666464484
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1666464484
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1666464484
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_227
timestamp 1666464484
transform 1 0 21988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1666464484
transform 1 0 22356 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1666464484
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_8
timestamp 1666464484
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1666464484
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1666464484
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1666464484
transform 1 0 22356 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_227
timestamp 1666464484
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1666464484
transform 1 0 22356 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1666464484
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1666464484
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_227
timestamp 1666464484
transform 1 0 21988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1666464484
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1666464484
transform 1 0 22356 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1666464484
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1666464484
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1666464484
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_231
timestamp 1666464484
transform 1 0 22356 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_227
timestamp 1666464484
transform 1 0 21988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1666464484
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1666464484
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1666464484
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_227
timestamp 1666464484
transform 1 0 21988 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_231
timestamp 1666464484
transform 1 0 22356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1666464484
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1666464484
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_32
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1666464484
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_231
timestamp 1666464484
transform 1 0 22356 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1666464484
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1666464484
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_231
timestamp 1666464484
transform 1 0 22356 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1666464484
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_231
timestamp 1666464484
transform 1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_8
timestamp 1666464484
transform 1 0 1840 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_20
timestamp 1666464484
transform 1 0 2944 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_32
timestamp 1666464484
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1666464484
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1666464484
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1666464484
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_231
timestamp 1666464484
transform 1 0 22356 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_8
timestamp 1666464484
transform 1 0 1840 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_231
timestamp 1666464484
transform 1 0 22356 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_14
timestamp 1666464484
transform 1 0 2392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1666464484
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_34
timestamp 1666464484
transform 1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_49
timestamp 1666464484
transform 1 0 5612 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_54
timestamp 1666464484
transform 1 0 6072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_57
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_68
timestamp 1666464484
transform 1 0 7360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_76
timestamp 1666464484
transform 1 0 8096 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1666464484
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_95
timestamp 1666464484
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1666464484
transform 1 0 11224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_113
timestamp 1666464484
transform 1 0 11500 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_122
timestamp 1666464484
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1666464484
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1666464484
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1666464484
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_181
timestamp 1666464484
transform 1 0 17756 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_203
timestamp 1666464484
transform 1 0 19780 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_215
timestamp 1666464484
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_225
timestamp 1666464484
transform 1 0 21804 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_230
timestamp 1666464484
transform 1 0 22264 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 22816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 22816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 22816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 22816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 22816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 22816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 22816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 22816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_2
timestamp 1666464484
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_3
timestamp 1666464484
transform 1 0 22080 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_4
timestamp 1666464484
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_5
timestamp 1666464484
transform 1 0 22080 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_6
timestamp 1666464484
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_7
timestamp 1666464484
transform 1 0 22080 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_8
timestamp 1666464484
transform 1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_9
timestamp 1666464484
transform 1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_10
timestamp 1666464484
transform 1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_11
timestamp 1666464484
transform 1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_12
timestamp 1666464484
transform 1 0 22080 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_13
timestamp 1666464484
transform 1 0 22080 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_14
timestamp 1666464484
transform 1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_15
timestamp 1666464484
transform 1 0 22080 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_16
timestamp 1666464484
transform -1 0 22264 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_17
timestamp 1666464484
transform -1 0 19780 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_18
timestamp 1666464484
transform -1 0 17756 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_19
timestamp 1666464484
transform -1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_20
timestamp 1666464484
transform -1 0 12328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_21
timestamp 1666464484
transform -1 0 9844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_22
timestamp 1666464484
transform -1 0 7360 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_23
timestamp 1666464484
transform -1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24
timestamp 1666464484
transform -1 0 2392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform -1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform -1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform -1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform -1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform 1 0 22080 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform 1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform 1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform 1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform 1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform 1 0 22080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform 1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform 1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform 1 0 22080 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform 1 0 22080 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform 1 0 22080 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform -1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform -1 0 18952 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform -1 0 17112 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform -1 0 14536 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform 1 0 10948 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform 1 0 8372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform 1 0 5796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform -1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform -1 0 1840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform -1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 23200 2864 24000 2984 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 23200 19184 24000 19304 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 23200 20816 24000 20936 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 23200 22448 24000 22568 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 23200 24080 24000 24200 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 23200 25712 24000 25832 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 22742 29200 22798 30000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 20258 29200 20314 30000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 17774 29200 17830 30000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 15290 29200 15346 30000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 12806 29200 12862 30000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 23200 4496 24000 4616 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 7838 29200 7894 30000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 5354 29200 5410 30000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 2870 29200 2926 30000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 23200 6128 24000 6248 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 23200 7760 24000 7880 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 23200 9392 24000 9512 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 23200 11024 24000 11144 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 23200 12656 24000 12776 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 23200 14288 24000 14408 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 23200 15920 24000 16040 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 23200 17552 24000 17672 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 23200 3952 24000 4072 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 23200 20272 24000 20392 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 23200 21904 24000 22024 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 23200 23536 24000 23656 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 23200 25168 24000 25288 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 23200 26800 24000 26920 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 21086 29200 21142 30000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 18602 29200 18658 30000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 13634 29200 13690 30000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 11150 29200 11206 30000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 23200 5584 24000 5704 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 8666 29200 8722 30000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 6182 29200 6238 30000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 3698 29200 3754 30000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 1214 29200 1270 30000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 23200 7216 24000 7336 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 23200 8848 24000 8968 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 23200 10480 24000 10600 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 23200 12112 24000 12232 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 23200 13744 24000 13864 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 23200 15376 24000 15496 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 23200 17008 24000 17128 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 23200 18640 24000 18760 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 23200 3408 24000 3528 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 23200 19728 24000 19848 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 23200 21360 24000 21480 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 23200 22992 24000 23112 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 23200 24624 24000 24744 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 23200 26256 24000 26376 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 19430 29200 19486 30000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 16946 29200 17002 30000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 14462 29200 14518 30000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 11978 29200 12034 30000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 23200 5040 24000 5160 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 9494 29200 9550 30000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 7010 29200 7066 30000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 2042 29200 2098 30000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 23200 6672 24000 6792 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 23200 8304 24000 8424 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 23200 9936 24000 10056 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 23200 11568 24000 11688 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 23200 13200 24000 13320 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 23200 14832 24000 14952 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 23200 16464 24000 16584 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 23200 18096 24000 18216 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 3658 2128 3978 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 9086 2128 9406 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 14514 2128 14834 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 19942 2128 20262 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 6372 2128 6692 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 11960 27744 11960 27744 0 vccd1
rlabel via1 12040 27200 12040 27200 0 vssd1
rlabel via2 22310 3485 22310 3485 0 net1
rlabel via2 22310 18139 22310 18139 0 net10
rlabel via2 22310 19805 22310 19805 0 net11
rlabel via2 22310 21403 22310 21403 0 net12
rlabel via2 22310 23069 22310 23069 0 net13
rlabel via2 22310 24667 22310 24667 0 net14
rlabel via2 22310 26333 22310 26333 0 net15
rlabel metal2 22034 28441 22034 28441 0 net16
rlabel metal2 19550 28441 19550 28441 0 net17
rlabel metal1 17250 27574 17250 27574 0 net18
rlabel metal2 14950 28441 14950 28441 0 net19
rlabel via2 22310 5083 22310 5083 0 net2
rlabel metal2 12098 28441 12098 28441 0 net20
rlabel metal2 9614 28441 9614 28441 0 net21
rlabel metal2 7130 28441 7130 28441 0 net22
rlabel metal2 4646 28441 4646 28441 0 net23
rlabel metal2 2162 28441 2162 28441 0 net24
rlabel metal1 2852 27574 2852 27574 0 net25
rlabel metal3 1142 26180 1142 26180 0 net26
rlabel metal3 1142 24140 1142 24140 0 net27
rlabel metal3 1142 22100 1142 22100 0 net28
rlabel metal3 1142 20060 1142 20060 0 net29
rlabel via2 22310 6749 22310 6749 0 net3
rlabel metal3 1142 18020 1142 18020 0 net30
rlabel metal3 1142 15980 1142 15980 0 net31
rlabel metal3 1142 13940 1142 13940 0 net32
rlabel metal3 1142 11900 1142 11900 0 net33
rlabel metal3 1142 9860 1142 9860 0 net34
rlabel metal3 1142 7820 1142 7820 0 net35
rlabel metal3 1142 5780 1142 5780 0 net36
rlabel metal3 1142 3740 1142 3740 0 net37
rlabel metal3 1142 1700 1142 1700 0 net38
rlabel via2 22310 3995 22310 3995 0 net39
rlabel via2 22310 8347 22310 8347 0 net4
rlabel via2 22310 5661 22310 5661 0 net40
rlabel via2 22310 7259 22310 7259 0 net41
rlabel via2 22310 8925 22310 8925 0 net42
rlabel via2 22310 10523 22310 10523 0 net43
rlabel via2 22310 12189 22310 12189 0 net44
rlabel via2 22310 13821 22310 13821 0 net45
rlabel via2 22310 15453 22310 15453 0 net46
rlabel via2 22310 17051 22310 17051 0 net47
rlabel via2 22310 18717 22310 18717 0 net48
rlabel via2 22310 20315 22310 20315 0 net49
rlabel via2 22310 10013 22310 10013 0 net5
rlabel metal2 22310 22049 22310 22049 0 net50
rlabel via2 22310 23579 22310 23579 0 net51
rlabel via2 22310 25245 22310 25245 0 net52
rlabel via2 22310 26843 22310 26843 0 net53
rlabel metal2 21206 28441 21206 28441 0 net54
rlabel metal2 18722 28441 18722 28441 0 net55
rlabel metal1 16744 27574 16744 27574 0 net56
rlabel metal1 14076 27574 14076 27574 0 net57
rlabel metal2 11178 28434 11178 28434 0 net58
rlabel metal2 8602 28441 8602 28441 0 net59
rlabel via2 22310 11611 22310 11611 0 net6
rlabel metal2 6026 28441 6026 28441 0 net60
rlabel metal1 4048 27574 4048 27574 0 net61
rlabel metal1 1518 26962 1518 26962 0 net62
rlabel metal1 2530 26962 2530 26962 0 net63
rlabel metal3 1142 25500 1142 25500 0 net64
rlabel metal3 1142 23460 1142 23460 0 net65
rlabel metal3 1142 21420 1142 21420 0 net66
rlabel metal3 1142 19380 1142 19380 0 net67
rlabel metal3 1142 17340 1142 17340 0 net68
rlabel metal3 1142 15300 1142 15300 0 net69
rlabel via2 22310 13277 22310 13277 0 net7
rlabel metal3 1142 13260 1142 13260 0 net70
rlabel metal3 1142 11220 1142 11220 0 net71
rlabel metal3 1142 9180 1142 9180 0 net72
rlabel metal3 1142 7140 1142 7140 0 net73
rlabel metal3 1142 5100 1142 5100 0 net74
rlabel metal3 1142 3060 1142 3060 0 net75
rlabel metal3 1050 1020 1050 1020 0 net76
rlabel via2 22310 14875 22310 14875 0 net8
rlabel metal2 22310 16575 22310 16575 0 net9
<< properties >>
string FIXED_BBOX 0 0 24000 30000
<< end >>
