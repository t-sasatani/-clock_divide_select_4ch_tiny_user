magic
tech sky130A
magscale 1 2
timestamp 1672368810
<< viali >>
rect 4997 17289 5031 17323
rect 10701 17289 10735 17323
rect 13093 17289 13127 17323
rect 5825 17221 5859 17255
rect 6653 17221 6687 17255
rect 1849 17153 1883 17187
rect 4445 17153 4479 17187
rect 6745 17153 6779 17187
rect 8329 17153 8363 17187
rect 9137 17153 9171 17187
rect 9505 17153 9539 17187
rect 10057 17153 10091 17187
rect 10977 17153 11011 17187
rect 11969 17153 12003 17187
rect 13737 17153 13771 17187
rect 15200 17153 15234 17187
rect 17224 17153 17258 17187
rect 1593 17085 1627 17119
rect 8585 17085 8619 17119
rect 10241 17085 10275 17119
rect 11713 17085 11747 17119
rect 14933 17085 14967 17119
rect 16957 17085 16991 17119
rect 5457 17017 5491 17051
rect 13553 17017 13587 17051
rect 2973 16949 3007 16983
rect 3985 16949 4019 16983
rect 4353 16949 4387 16983
rect 5825 16949 5859 16983
rect 6009 16949 6043 16983
rect 7205 16949 7239 16983
rect 14289 16949 14323 16983
rect 16313 16949 16347 16983
rect 18337 16949 18371 16983
rect 6561 16745 6595 16779
rect 12357 16745 12391 16779
rect 5089 16677 5123 16711
rect 6745 16677 6779 16711
rect 13001 16677 13035 16711
rect 2973 16609 3007 16643
rect 6193 16609 6227 16643
rect 16773 16609 16807 16643
rect 17325 16609 17359 16643
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 4353 16541 4387 16575
rect 5457 16541 5491 16575
rect 7205 16541 7239 16575
rect 10517 16541 10551 16575
rect 10977 16541 11011 16575
rect 16037 16541 16071 16575
rect 17049 16541 17083 16575
rect 17417 16541 17451 16575
rect 17785 16541 17819 16575
rect 18337 16541 18371 16575
rect 2728 16473 2762 16507
rect 4261 16473 4295 16507
rect 6561 16473 6595 16507
rect 7472 16473 7506 16507
rect 10250 16473 10284 16507
rect 11244 16473 11278 16507
rect 13277 16473 13311 16507
rect 15792 16473 15826 16507
rect 1593 16405 1627 16439
rect 4537 16405 4571 16439
rect 4997 16405 5031 16439
rect 8585 16405 8619 16439
rect 9137 16405 9171 16439
rect 12817 16405 12851 16439
rect 14657 16405 14691 16439
rect 2973 16201 3007 16235
rect 4997 16201 5031 16235
rect 10149 16201 10183 16235
rect 12633 16201 12667 16235
rect 16313 16201 16347 16235
rect 18337 16201 18371 16235
rect 4813 16133 4847 16167
rect 7113 16133 7147 16167
rect 7941 16133 7975 16167
rect 8029 16133 8063 16167
rect 14105 16133 14139 16167
rect 14197 16133 14231 16167
rect 15178 16133 15212 16167
rect 17202 16133 17236 16167
rect 1593 16065 1627 16099
rect 1860 16065 1894 16099
rect 3617 16065 3651 16099
rect 3709 16065 3743 16099
rect 3985 16065 4019 16099
rect 7777 16065 7811 16099
rect 8171 16065 8205 16099
rect 8769 16065 8803 16099
rect 9036 16065 9070 16099
rect 10793 16065 10827 16099
rect 10885 16065 10919 16099
rect 11161 16065 11195 16099
rect 12817 16065 12851 16099
rect 13001 16065 13035 16099
rect 13093 16065 13127 16099
rect 13921 16065 13955 16099
rect 14289 16065 14323 16099
rect 16957 16065 16991 16099
rect 5457 15997 5491 16031
rect 5917 15997 5951 16031
rect 11069 15997 11103 16031
rect 12173 15997 12207 16031
rect 14933 15997 14967 16031
rect 4445 15929 4479 15963
rect 5641 15929 5675 15963
rect 6745 15929 6779 15963
rect 11805 15929 11839 15963
rect 3433 15861 3467 15895
rect 3893 15861 3927 15895
rect 4813 15861 4847 15895
rect 7113 15861 7147 15895
rect 7297 15861 7331 15895
rect 8309 15861 8343 15895
rect 10609 15861 10643 15895
rect 11713 15861 11747 15895
rect 14473 15861 14507 15895
rect 11253 15657 11287 15691
rect 12909 15657 12943 15691
rect 14289 15657 14323 15691
rect 15025 15657 15059 15691
rect 15485 15657 15519 15691
rect 16313 15657 16347 15691
rect 7389 15589 7423 15623
rect 11897 15589 11931 15623
rect 13553 15589 13587 15623
rect 18337 15589 18371 15623
rect 2421 15521 2455 15555
rect 3985 15521 4019 15555
rect 8125 15521 8159 15555
rect 1593 15453 1627 15487
rect 2513 15453 2547 15487
rect 2973 15453 3007 15487
rect 3433 15453 3467 15487
rect 4241 15453 4275 15487
rect 5825 15453 5859 15487
rect 6101 15453 6135 15487
rect 8033 15453 8067 15487
rect 8308 15453 8342 15487
rect 8401 15453 8435 15487
rect 8585 15453 8619 15487
rect 10517 15453 10551 15487
rect 11437 15453 11471 15487
rect 14473 15453 14507 15487
rect 14933 15453 14967 15487
rect 15209 15453 15243 15487
rect 15301 15453 15335 15487
rect 15945 15453 15979 15487
rect 16957 15453 16991 15487
rect 6285 15385 6319 15419
rect 7113 15385 7147 15419
rect 10272 15385 10306 15419
rect 12081 15385 12115 15419
rect 12265 15385 12299 15419
rect 12877 15385 12911 15419
rect 13093 15385 13127 15419
rect 16313 15385 16347 15419
rect 17224 15385 17258 15419
rect 1869 15317 1903 15351
rect 5365 15317 5399 15351
rect 5917 15317 5951 15351
rect 7573 15317 7607 15351
rect 9137 15317 9171 15351
rect 10977 15317 11011 15351
rect 12725 15317 12759 15351
rect 16497 15317 16531 15351
rect 2973 15113 3007 15147
rect 5089 15113 5123 15147
rect 9781 15113 9815 15147
rect 18337 15113 18371 15147
rect 5549 15045 5583 15079
rect 5765 15045 5799 15079
rect 6837 15045 6871 15079
rect 7817 15045 7851 15079
rect 8033 15045 8067 15079
rect 10149 15045 10183 15079
rect 11881 15045 11915 15079
rect 12081 15045 12115 15079
rect 13369 15045 13403 15079
rect 14181 15045 14215 15079
rect 14355 15045 14389 15079
rect 17202 15045 17236 15079
rect 1593 14977 1627 15011
rect 1860 14977 1894 15011
rect 3612 14977 3646 15011
rect 3709 14977 3743 15011
rect 3801 14977 3835 15011
rect 3984 14977 4018 15011
rect 4077 14977 4111 15011
rect 4537 14977 4571 15011
rect 4813 14977 4847 15011
rect 4905 14977 4939 15011
rect 7021 14977 7055 15011
rect 8861 14977 8895 15011
rect 9960 14977 9994 15011
rect 10057 14977 10091 15011
rect 10332 14977 10366 15011
rect 10425 14977 10459 15011
rect 11161 14977 11195 15011
rect 12541 14977 12575 15011
rect 13553 14977 13587 15011
rect 15761 14977 15795 15011
rect 16037 14977 16071 15011
rect 16129 14977 16163 15011
rect 8769 14909 8803 14943
rect 14841 14909 14875 14943
rect 16957 14909 16991 14943
rect 3433 14841 3467 14875
rect 7205 14841 7239 14875
rect 14013 14841 14047 14875
rect 15209 14841 15243 14875
rect 15301 14841 15335 14875
rect 4629 14773 4663 14807
rect 5733 14773 5767 14807
rect 5917 14773 5951 14807
rect 7665 14773 7699 14807
rect 7849 14773 7883 14807
rect 8585 14773 8619 14807
rect 10977 14773 11011 14807
rect 11713 14773 11747 14807
rect 11897 14773 11931 14807
rect 13185 14773 13219 14807
rect 14197 14773 14231 14807
rect 15853 14773 15887 14807
rect 16313 14773 16347 14807
rect 4169 14569 4203 14603
rect 5825 14569 5859 14603
rect 6837 14569 6871 14603
rect 8401 14569 8435 14603
rect 9321 14569 9355 14603
rect 12449 14569 12483 14603
rect 14289 14569 14323 14603
rect 15853 14569 15887 14603
rect 16865 14569 16899 14603
rect 3985 14501 4019 14535
rect 17233 14501 17267 14535
rect 6193 14433 6227 14467
rect 11989 14433 12023 14467
rect 16221 14433 16255 14467
rect 1593 14365 1627 14399
rect 4537 14365 4571 14399
rect 6009 14365 6043 14399
rect 6768 14365 6802 14399
rect 6929 14365 6963 14399
rect 7573 14365 7607 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 13093 14365 13127 14399
rect 14933 14365 14967 14399
rect 15761 14365 15795 14399
rect 17831 14365 17865 14399
rect 18061 14365 18095 14399
rect 18244 14365 18278 14399
rect 18337 14365 18371 14399
rect 1860 14297 1894 14331
rect 5181 14297 5215 14331
rect 5365 14297 5399 14331
rect 7757 14297 7791 14331
rect 8217 14297 8251 14331
rect 8433 14297 8467 14331
rect 11722 14297 11756 14331
rect 13185 14297 13219 14331
rect 15117 14297 15151 14331
rect 15301 14297 15335 14331
rect 17969 14297 18003 14331
rect 2973 14229 3007 14263
rect 4169 14229 4203 14263
rect 4997 14229 5031 14263
rect 7389 14229 7423 14263
rect 8585 14229 8619 14263
rect 9689 14229 9723 14263
rect 10609 14229 10643 14263
rect 16681 14229 16715 14263
rect 16865 14229 16899 14263
rect 17693 14229 17727 14263
rect 2973 14025 3007 14059
rect 3893 14025 3927 14059
rect 4721 14025 4755 14059
rect 9873 14025 9907 14059
rect 10333 14025 10367 14059
rect 11713 14025 11747 14059
rect 15945 14025 15979 14059
rect 17785 14025 17819 14059
rect 4353 13957 4387 13991
rect 4569 13957 4603 13991
rect 6806 13957 6840 13991
rect 8738 13957 8772 13991
rect 10485 13957 10519 13991
rect 10701 13957 10735 13991
rect 15117 13957 15151 13991
rect 15333 13957 15367 13991
rect 16113 13957 16147 13991
rect 16313 13957 16347 13991
rect 17325 13957 17359 13991
rect 17969 13957 18003 13991
rect 1593 13889 1627 13923
rect 1860 13889 1894 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 3709 13889 3743 13923
rect 5535 13889 5569 13923
rect 12081 13889 12115 13923
rect 13369 13889 13403 13923
rect 14473 13889 14507 13923
rect 5457 13821 5491 13855
rect 6561 13821 6595 13855
rect 8493 13821 8527 13855
rect 12173 13821 12207 13855
rect 14013 13821 14047 13855
rect 16865 13821 16899 13855
rect 5825 13753 5859 13787
rect 15485 13753 15519 13787
rect 16957 13753 16991 13787
rect 18337 13753 18371 13787
rect 4537 13685 4571 13719
rect 7941 13685 7975 13719
rect 10517 13685 10551 13719
rect 15301 13685 15335 13719
rect 16129 13685 16163 13719
rect 17969 13685 18003 13719
rect 1961 13481 1995 13515
rect 4169 13481 4203 13515
rect 4353 13481 4387 13515
rect 5825 13481 5859 13515
rect 6009 13481 6043 13515
rect 6653 13481 6687 13515
rect 14657 13481 14691 13515
rect 15301 13481 15335 13515
rect 17417 13481 17451 13515
rect 18337 13481 18371 13515
rect 2145 13413 2179 13447
rect 2697 13413 2731 13447
rect 4813 13413 4847 13447
rect 8585 13413 8619 13447
rect 18153 13413 18187 13447
rect 3065 13345 3099 13379
rect 10231 13345 10265 13379
rect 10517 13345 10551 13379
rect 10793 13345 10827 13379
rect 13737 13345 13771 13379
rect 16497 13345 16531 13379
rect 1593 13277 1627 13311
rect 5181 13277 5215 13311
rect 7757 13277 7791 13311
rect 8401 13277 8435 13311
rect 10379 13277 10413 13311
rect 11253 13277 11287 13311
rect 11437 13277 11471 13311
rect 11897 13277 11931 13311
rect 12909 13277 12943 13311
rect 14841 13277 14875 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 16957 13277 16991 13311
rect 17049 13277 17083 13311
rect 17233 13277 17267 13311
rect 3985 13209 4019 13243
rect 4997 13209 5031 13243
rect 5641 13209 5675 13243
rect 6469 13209 6503 13243
rect 8217 13209 8251 13243
rect 17877 13209 17911 13243
rect 1961 13141 1995 13175
rect 2605 13141 2639 13175
rect 4195 13141 4229 13175
rect 5841 13141 5875 13175
rect 6669 13141 6703 13175
rect 6837 13141 6871 13175
rect 7573 13141 7607 13175
rect 9597 13141 9631 13175
rect 13093 13141 13127 13175
rect 2145 12937 2179 12971
rect 4721 12937 4755 12971
rect 7941 12937 7975 12971
rect 8861 12937 8895 12971
rect 10333 12937 10367 12971
rect 10977 12937 11011 12971
rect 11805 12937 11839 12971
rect 13001 12937 13035 12971
rect 13737 12937 13771 12971
rect 17207 12937 17241 12971
rect 17877 12937 17911 12971
rect 18245 12937 18279 12971
rect 1961 12869 1995 12903
rect 4371 12869 4405 12903
rect 4537 12869 4571 12903
rect 6806 12869 6840 12903
rect 17417 12869 17451 12903
rect 1593 12801 1627 12835
rect 3709 12801 3743 12835
rect 5641 12801 5675 12835
rect 9045 12801 9079 12835
rect 9137 12801 9171 12835
rect 9873 12801 9907 12835
rect 10517 12801 10551 12835
rect 11161 12801 11195 12835
rect 12265 12801 12299 12835
rect 13093 12801 13127 12835
rect 13553 12801 13587 12835
rect 13737 12801 13771 12835
rect 14197 12801 14231 12835
rect 15025 12801 15059 12835
rect 15669 12801 15703 12835
rect 18061 12801 18095 12835
rect 18337 12801 18371 12835
rect 2605 12733 2639 12767
rect 3065 12733 3099 12767
rect 3525 12733 3559 12767
rect 5549 12733 5583 12767
rect 6561 12733 6595 12767
rect 2973 12665 3007 12699
rect 6009 12665 6043 12699
rect 12449 12665 12483 12699
rect 15485 12665 15519 12699
rect 16313 12665 16347 12699
rect 1961 12597 1995 12631
rect 3893 12597 3927 12631
rect 9689 12597 9723 12631
rect 14381 12597 14415 12631
rect 17049 12597 17083 12631
rect 17233 12597 17267 12631
rect 4997 12393 5031 12427
rect 6561 12393 6595 12427
rect 7205 12393 7239 12427
rect 9229 12393 9263 12427
rect 9873 12393 9907 12427
rect 10701 12393 10735 12427
rect 11805 12393 11839 12427
rect 14749 12393 14783 12427
rect 16681 12393 16715 12427
rect 17233 12393 17267 12427
rect 18061 12393 18095 12427
rect 6009 12325 6043 12359
rect 13737 12325 13771 12359
rect 15393 12325 15427 12359
rect 1593 12257 1627 12291
rect 16037 12257 16071 12291
rect 3985 12189 4019 12223
rect 5641 12189 5675 12223
rect 6653 12189 6687 12223
rect 7113 12189 7147 12223
rect 7757 12189 7791 12223
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 9413 12189 9447 12223
rect 10057 12189 10091 12223
rect 10517 12189 10551 12223
rect 11161 12189 11195 12223
rect 11989 12189 12023 12223
rect 13093 12189 13127 12223
rect 14565 12189 14599 12223
rect 15209 12189 15243 12223
rect 1860 12121 1894 12155
rect 4169 12121 4203 12155
rect 4353 12121 4387 12155
rect 4981 12121 5015 12155
rect 5181 12121 5215 12155
rect 5825 12121 5859 12155
rect 17325 12121 17359 12155
rect 18029 12121 18063 12155
rect 18245 12121 18279 12155
rect 2973 12053 3007 12087
rect 4813 12053 4847 12087
rect 7941 12053 7975 12087
rect 8585 12053 8619 12087
rect 17877 12053 17911 12087
rect 6653 11849 6687 11883
rect 9137 11849 9171 11883
rect 9597 11849 9631 11883
rect 10333 11849 10367 11883
rect 10885 11849 10919 11883
rect 14289 11849 14323 11883
rect 14933 11849 14967 11883
rect 15669 11849 15703 11883
rect 17969 11849 18003 11883
rect 5533 11781 5567 11815
rect 5733 11781 5767 11815
rect 18337 11781 18371 11815
rect 1593 11713 1627 11747
rect 1860 11713 1894 11747
rect 3433 11713 3467 11747
rect 3709 11713 3743 11747
rect 3801 11713 3835 11747
rect 4905 11713 4939 11747
rect 7113 11713 7147 11747
rect 7849 11713 7883 11747
rect 8953 11713 8987 11747
rect 9781 11713 9815 11747
rect 10241 11713 10275 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 13737 11713 13771 11747
rect 14381 11713 14415 11747
rect 14841 11713 14875 11747
rect 15485 11713 15519 11747
rect 15669 11713 15703 11747
rect 16313 11713 16347 11747
rect 18153 11713 18187 11747
rect 3525 11645 3559 11679
rect 3985 11645 4019 11679
rect 13093 11645 13127 11679
rect 5365 11577 5399 11611
rect 17509 11577 17543 11611
rect 2973 11509 3007 11543
rect 4445 11509 4479 11543
rect 4629 11509 4663 11543
rect 5549 11509 5583 11543
rect 3985 11305 4019 11339
rect 4169 11305 4203 11339
rect 6837 11305 6871 11339
rect 7297 11305 7331 11339
rect 9137 11305 9171 11339
rect 9781 11305 9815 11339
rect 13645 11305 13679 11339
rect 15117 11305 15151 11339
rect 16221 11305 16255 11339
rect 17049 11305 17083 11339
rect 17509 11305 17543 11339
rect 2973 11237 3007 11271
rect 7941 11237 7975 11271
rect 11069 11237 11103 11271
rect 14473 11237 14507 11271
rect 15669 11237 15703 11271
rect 1593 11169 1627 11203
rect 10425 11169 10459 11203
rect 4537 11101 4571 11135
rect 4997 11101 5031 11135
rect 5273 11101 5307 11135
rect 6101 11101 6135 11135
rect 6653 11101 6687 11135
rect 8125 11101 8159 11135
rect 9321 11101 9355 11135
rect 9965 11101 9999 11135
rect 15761 11101 15795 11135
rect 16405 11101 16439 11135
rect 16865 11101 16899 11135
rect 17693 11101 17727 11135
rect 18337 11101 18371 11135
rect 1860 11033 1894 11067
rect 5457 11033 5491 11067
rect 5917 11033 5951 11067
rect 11713 11033 11747 11067
rect 4169 10965 4203 10999
rect 5089 10965 5123 10999
rect 18153 10965 18187 10999
rect 6929 10761 6963 10795
rect 9321 10761 9355 10795
rect 10057 10761 10091 10795
rect 15025 10761 15059 10795
rect 17509 10761 17543 10795
rect 2145 10625 2179 10659
rect 2513 10625 2547 10659
rect 2881 10625 2915 10659
rect 3433 10625 3467 10659
rect 5017 10625 5051 10659
rect 5273 10625 5307 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 6745 10625 6779 10659
rect 7389 10625 7423 10659
rect 8677 10625 8711 10659
rect 9505 10625 9539 10659
rect 9965 10625 9999 10659
rect 15669 10625 15703 10659
rect 16865 10625 16899 10659
rect 17693 10625 17727 10659
rect 18337 10625 18371 10659
rect 2053 10557 2087 10591
rect 2421 10557 2455 10591
rect 8033 10557 8067 10591
rect 10609 10557 10643 10591
rect 16313 10557 16347 10591
rect 3893 10489 3927 10523
rect 17049 10489 17083 10523
rect 5733 10421 5767 10455
rect 4629 10217 4663 10251
rect 5457 10217 5491 10251
rect 6745 10217 6779 10251
rect 8125 10217 8159 10251
rect 9137 10217 9171 10251
rect 9781 10217 9815 10251
rect 15669 10217 15703 10251
rect 16313 10217 16347 10251
rect 17417 10217 17451 10251
rect 18337 10217 18371 10251
rect 16773 10149 16807 10183
rect 1593 10081 1627 10115
rect 7481 10081 7515 10115
rect 3985 10013 4019 10047
rect 4078 10013 4112 10047
rect 4261 10013 4295 10047
rect 4491 10013 4525 10047
rect 5273 10013 5307 10047
rect 6285 10013 6319 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 8033 10013 8067 10047
rect 9321 10013 9355 10047
rect 16957 10013 16991 10047
rect 17601 10013 17635 10047
rect 1860 9945 1894 9979
rect 4353 9945 4387 9979
rect 5089 9945 5123 9979
rect 2973 9877 3007 9911
rect 6101 9877 6135 9911
rect 7849 9673 7883 9707
rect 3709 9605 3743 9639
rect 4905 9605 4939 9639
rect 5733 9605 5767 9639
rect 9781 9605 9815 9639
rect 16313 9605 16347 9639
rect 1593 9537 1627 9571
rect 1860 9537 1894 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 3801 9537 3835 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 6745 9537 6779 9571
rect 8033 9537 8067 9571
rect 8677 9537 8711 9571
rect 9137 9537 9171 9571
rect 15761 9537 15795 9571
rect 17049 9537 17083 9571
rect 17693 9537 17727 9571
rect 18337 9537 18371 9571
rect 4445 9469 4479 9503
rect 2973 9401 3007 9435
rect 3985 9401 4019 9435
rect 4629 9401 4663 9435
rect 7205 9401 7239 9435
rect 16865 9401 16899 9435
rect 17509 9401 17543 9435
rect 6561 9333 6595 9367
rect 8493 9333 8527 9367
rect 5549 9129 5583 9163
rect 6837 9129 6871 9163
rect 7481 9129 7515 9163
rect 8125 9129 8159 9163
rect 9137 9129 9171 9163
rect 17141 9129 17175 9163
rect 18337 9129 18371 9163
rect 4077 9061 4111 9095
rect 4905 9061 4939 9095
rect 6377 9061 6411 9095
rect 16681 9061 16715 9095
rect 16129 8993 16163 9027
rect 2973 8925 3007 8959
rect 6193 8925 6227 8959
rect 7021 8925 7055 8959
rect 2728 8857 2762 8891
rect 4445 8857 4479 8891
rect 1593 8789 1627 8823
rect 3985 8789 4019 8823
rect 2145 8585 2179 8619
rect 2973 8585 3007 8619
rect 3893 8585 3927 8619
rect 4537 8585 4571 8619
rect 17325 8585 17359 8619
rect 1961 8517 1995 8551
rect 3525 8517 3559 8551
rect 3730 8517 3764 8551
rect 1593 8449 1627 8483
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 4353 8449 4387 8483
rect 4997 8449 5031 8483
rect 5825 8449 5859 8483
rect 6745 8449 6779 8483
rect 7205 8449 7239 8483
rect 18337 8449 18371 8483
rect 7849 8381 7883 8415
rect 2605 8313 2639 8347
rect 6561 8313 6595 8347
rect 1961 8245 1995 8279
rect 3709 8245 3743 8279
rect 5181 8245 5215 8279
rect 5641 8245 5675 8279
rect 1593 8041 1627 8075
rect 2053 8041 2087 8075
rect 2605 8041 2639 8075
rect 2789 8041 2823 8075
rect 3985 8041 4019 8075
rect 4721 8041 4755 8075
rect 5273 8041 5307 8075
rect 6745 8041 6779 8075
rect 7205 7973 7239 8007
rect 18337 7905 18371 7939
rect 1777 7837 1811 7871
rect 1869 7837 1903 7871
rect 2145 7837 2179 7871
rect 4813 7837 4847 7871
rect 5917 7837 5951 7871
rect 6561 7837 6595 7871
rect 2773 7769 2807 7803
rect 2973 7769 3007 7803
rect 2421 7497 2455 7531
rect 3065 7497 3099 7531
rect 5641 7497 5675 7531
rect 6561 7497 6595 7531
rect 7113 7497 7147 7531
rect 1593 7429 1627 7463
rect 1809 7429 1843 7463
rect 2605 7361 2639 7395
rect 3249 7361 3283 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 5825 7361 5859 7395
rect 18337 7361 18371 7395
rect 3709 7293 3743 7327
rect 4997 7293 5031 7327
rect 1961 7225 1995 7259
rect 1777 7157 1811 7191
rect 4445 7157 4479 7191
rect 6009 6953 6043 6987
rect 4629 6885 4663 6919
rect 4077 6817 4111 6851
rect 1593 6749 1627 6783
rect 2421 6749 2455 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 4169 6749 4203 6783
rect 4813 6749 4847 6783
rect 5549 6749 5583 6783
rect 18337 6749 18371 6783
rect 1777 6613 1811 6647
rect 2237 6613 2271 6647
rect 3065 6613 3099 6647
rect 1777 6409 1811 6443
rect 3617 6409 3651 6443
rect 4813 6409 4847 6443
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 2881 6273 2915 6307
rect 3709 6273 3743 6307
rect 4353 6273 4387 6307
rect 5365 6273 5399 6307
rect 18337 6273 18371 6307
rect 2421 6137 2455 6171
rect 4169 6137 4203 6171
rect 2237 5865 2271 5899
rect 2881 5865 2915 5899
rect 4629 5865 4663 5899
rect 1685 5797 1719 5831
rect 1777 5661 1811 5695
rect 2421 5661 2455 5695
rect 3985 5661 4019 5695
rect 18337 5661 18371 5695
rect 1685 5321 1719 5355
rect 1777 5185 1811 5219
rect 2237 5185 2271 5219
rect 2881 5185 2915 5219
rect 18337 5049 18371 5083
rect 1869 4573 1903 4607
rect 18337 4573 18371 4607
rect 1685 4437 1719 4471
rect 1593 4097 1627 4131
rect 18337 3893 18371 3927
rect 1593 3689 1627 3723
rect 18337 3485 18371 3519
rect 1593 3009 1627 3043
rect 18337 2805 18371 2839
rect 1593 2601 1627 2635
rect 2237 2397 2271 2431
rect 2881 2397 2915 2431
rect 17693 2397 17727 2431
rect 18337 2397 18371 2431
<< metal1 >>
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 13538 17728 13544 17740
rect 10008 17700 13544 17728
rect 10008 17688 10014 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 10502 17660 10508 17672
rect 8628 17632 10508 17660
rect 8628 17620 8634 17632
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 6546 17552 6552 17604
rect 6604 17592 6610 17604
rect 10594 17592 10600 17604
rect 6604 17564 10600 17592
rect 6604 17552 6610 17564
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 7098 17524 7104 17536
rect 5592 17496 7104 17524
rect 5592 17484 5598 17496
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10686 17524 10692 17536
rect 9732 17496 10692 17524
rect 9732 17484 9738 17496
rect 10686 17484 10692 17496
rect 10744 17524 10750 17536
rect 13722 17524 13728 17536
rect 10744 17496 13728 17524
rect 10744 17484 10750 17496
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 18782 17484 18788 17536
rect 18840 17524 18846 17536
rect 19426 17524 19432 17536
rect 18840 17496 19432 17524
rect 18840 17484 18846 17496
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 9674 17320 9680 17332
rect 5031 17292 9680 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10594 17280 10600 17332
rect 10652 17320 10658 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10652 17292 10701 17320
rect 10652 17280 10658 17292
rect 10689 17289 10701 17292
rect 10735 17320 10747 17323
rect 11238 17320 11244 17332
rect 10735 17292 11244 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 12406 17292 13093 17320
rect 5813 17255 5871 17261
rect 5813 17221 5825 17255
rect 5859 17252 5871 17255
rect 6546 17252 6552 17264
rect 5859 17224 6552 17252
rect 5859 17221 5871 17224
rect 5813 17215 5871 17221
rect 6546 17212 6552 17224
rect 6604 17212 6610 17264
rect 6641 17255 6699 17261
rect 6641 17221 6653 17255
rect 6687 17252 6699 17255
rect 10778 17252 10784 17264
rect 6687 17224 10784 17252
rect 6687 17221 6699 17224
rect 6641 17215 6699 17221
rect 10778 17212 10784 17224
rect 10836 17212 10842 17264
rect 12406 17252 12434 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13081 17283 13139 17289
rect 10980 17224 12434 17252
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1837 17187 1895 17193
rect 1837 17184 1849 17187
rect 992 17156 1849 17184
rect 992 17144 998 17156
rect 1837 17153 1849 17156
rect 1883 17153 1895 17187
rect 1837 17147 1895 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 5718 17184 5724 17196
rect 4479 17156 5724 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 8317 17187 8375 17193
rect 8317 17153 8329 17187
rect 8363 17184 8375 17187
rect 9122 17184 9128 17196
rect 8363 17156 8708 17184
rect 9083 17156 9128 17184
rect 8363 17153 8375 17156
rect 8317 17147 8375 17153
rect 1486 17076 1492 17128
rect 1544 17116 1550 17128
rect 1581 17119 1639 17125
rect 1581 17116 1593 17119
rect 1544 17088 1593 17116
rect 1544 17076 1550 17088
rect 1581 17085 1593 17088
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 3016 17088 6684 17116
rect 3016 17076 3022 17088
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 5445 17051 5503 17057
rect 5445 17048 5457 17051
rect 5132 17020 5457 17048
rect 5132 17008 5138 17020
rect 5445 17017 5457 17020
rect 5491 17017 5503 17051
rect 5445 17011 5503 17017
rect 2961 16983 3019 16989
rect 2961 16949 2973 16983
rect 3007 16980 3019 16983
rect 3510 16980 3516 16992
rect 3007 16952 3516 16980
rect 3007 16949 3019 16952
rect 2961 16943 3019 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 3973 16983 4031 16989
rect 3973 16980 3985 16983
rect 3844 16952 3985 16980
rect 3844 16940 3850 16952
rect 3973 16949 3985 16952
rect 4019 16949 4031 16983
rect 3973 16943 4031 16949
rect 4341 16983 4399 16989
rect 4341 16949 4353 16983
rect 4387 16980 4399 16983
rect 5166 16980 5172 16992
rect 4387 16952 5172 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5813 16983 5871 16989
rect 5813 16949 5825 16983
rect 5859 16980 5871 16983
rect 5902 16980 5908 16992
rect 5859 16952 5908 16980
rect 5859 16949 5871 16952
rect 5813 16943 5871 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6656 16980 6684 17088
rect 6748 17048 6776 17147
rect 8570 17116 8576 17128
rect 8531 17088 8576 17116
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8680 17048 8708 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 9364 17156 9505 17184
rect 9364 17144 9370 17156
rect 9493 17153 9505 17156
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10980 17193 11008 17224
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 9732 17156 10057 17184
rect 9732 17144 9738 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11957 17187 12015 17193
rect 11957 17184 11969 17187
rect 11112 17156 11969 17184
rect 11112 17144 11118 17156
rect 11957 17153 11969 17156
rect 12003 17153 12015 17187
rect 13722 17184 13728 17196
rect 13683 17156 13728 17184
rect 11957 17147 12015 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 15194 17193 15200 17196
rect 15188 17147 15200 17193
rect 15252 17184 15258 17196
rect 17212 17187 17270 17193
rect 15252 17156 15288 17184
rect 15194 17144 15200 17147
rect 15252 17144 15258 17156
rect 17212 17153 17224 17187
rect 17258 17184 17270 17187
rect 17954 17184 17960 17196
rect 17258 17156 17960 17184
rect 17258 17153 17270 17156
rect 17212 17147 17270 17153
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 10229 17119 10287 17125
rect 10229 17085 10241 17119
rect 10275 17116 10287 17119
rect 10318 17116 10324 17128
rect 10275 17088 10324 17116
rect 10275 17085 10287 17088
rect 10229 17079 10287 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 10560 17088 11713 17116
rect 10560 17076 10566 17088
rect 11701 17085 11713 17088
rect 11747 17085 11759 17119
rect 14918 17116 14924 17128
rect 14879 17088 14924 17116
rect 11701 17079 11759 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 16942 17116 16948 17128
rect 16903 17088 16948 17116
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 10410 17048 10416 17060
rect 6748 17020 7696 17048
rect 8680 17020 10416 17048
rect 6822 16980 6828 16992
rect 6052 16952 6097 16980
rect 6656 16952 6828 16980
rect 6052 16940 6058 16952
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7190 16980 7196 16992
rect 7151 16952 7196 16980
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 7668 16980 7696 17020
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 13541 17051 13599 17057
rect 13541 17048 13553 17051
rect 13004 17020 13553 17048
rect 13004 16980 13032 17020
rect 13541 17017 13553 17020
rect 13587 17017 13599 17051
rect 13541 17011 13599 17017
rect 14274 16980 14280 16992
rect 7668 16952 13032 16980
rect 14235 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 16298 16980 16304 16992
rect 16259 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 17184 16952 18337 16980
rect 17184 16940 17190 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 11146 16776 11152 16788
rect 6595 16748 11152 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 12342 16776 12348 16788
rect 11664 16748 11928 16776
rect 12255 16748 12348 16776
rect 11664 16736 11670 16748
rect 3510 16668 3516 16720
rect 3568 16708 3574 16720
rect 5077 16711 5135 16717
rect 5077 16708 5089 16711
rect 3568 16680 5089 16708
rect 3568 16668 3574 16680
rect 5077 16677 5089 16680
rect 5123 16677 5135 16711
rect 5077 16671 5135 16677
rect 6733 16711 6791 16717
rect 6733 16677 6745 16711
rect 6779 16677 6791 16711
rect 11900 16708 11928 16748
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 12618 16776 12624 16788
rect 12400 16748 12624 16776
rect 12400 16736 12406 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 15838 16776 15844 16788
rect 15028 16748 15844 16776
rect 12989 16711 13047 16717
rect 11900 16680 12434 16708
rect 6733 16671 6791 16677
rect 2958 16640 2964 16652
rect 2884 16612 2964 16640
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2884 16572 2912 16612
rect 2958 16600 2964 16612
rect 3016 16640 3022 16652
rect 6181 16643 6239 16649
rect 3016 16612 3109 16640
rect 4356 16612 5304 16640
rect 3016 16600 3022 16612
rect 4356 16584 4384 16612
rect 1728 16544 2912 16572
rect 1728 16532 1734 16544
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3936 16544 3985 16572
rect 3936 16532 3942 16544
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 3973 16535 4031 16541
rect 4081 16544 4169 16572
rect 2716 16507 2774 16513
rect 2716 16473 2728 16507
rect 2762 16504 2774 16507
rect 3326 16504 3332 16516
rect 2762 16476 3332 16504
rect 2762 16473 2774 16476
rect 2716 16467 2774 16473
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 4081 16436 4109 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4396 16544 4489 16572
rect 4396 16532 4402 16544
rect 4246 16504 4252 16516
rect 4207 16476 4252 16504
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 5276 16504 5304 16612
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6638 16640 6644 16652
rect 6227 16612 6644 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 6748 16640 6776 16671
rect 12406 16640 12434 16680
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 13078 16708 13084 16720
rect 13035 16680 13084 16708
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 13078 16668 13084 16680
rect 13136 16668 13142 16720
rect 15028 16640 15056 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 6748 16612 7328 16640
rect 12406 16612 15056 16640
rect 15948 16612 16773 16640
rect 7300 16584 7328 16612
rect 5442 16572 5448 16584
rect 5403 16544 5448 16572
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6822 16532 6828 16584
rect 6880 16572 6886 16584
rect 7193 16575 7251 16581
rect 7193 16572 7205 16575
rect 6880 16544 7205 16572
rect 6880 16532 6886 16544
rect 7193 16541 7205 16544
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 6178 16504 6184 16516
rect 5276 16476 6184 16504
rect 6178 16464 6184 16476
rect 6236 16464 6242 16516
rect 6546 16504 6552 16516
rect 6507 16476 6552 16504
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 7208 16504 7236 16535
rect 7282 16532 7288 16584
rect 7340 16532 7346 16584
rect 7392 16544 7880 16572
rect 7392 16504 7420 16544
rect 7208 16476 7420 16504
rect 7460 16507 7518 16513
rect 7460 16473 7472 16507
rect 7506 16473 7518 16507
rect 7852 16504 7880 16544
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 8996 16544 10364 16572
rect 8996 16532 9002 16544
rect 8662 16504 8668 16516
rect 7852 16476 8668 16504
rect 7460 16467 7518 16473
rect 4430 16436 4436 16448
rect 4081 16408 4436 16436
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 4890 16436 4896 16448
rect 4571 16408 4896 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5040 16408 5085 16436
rect 5040 16396 5046 16408
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7475 16436 7503 16467
rect 8662 16464 8668 16476
rect 8720 16464 8726 16516
rect 10226 16504 10232 16516
rect 10284 16513 10290 16516
rect 10196 16476 10232 16504
rect 10226 16464 10232 16476
rect 10284 16467 10296 16513
rect 10336 16504 10364 16544
rect 10502 16532 10508 16584
rect 10560 16572 10566 16584
rect 10686 16572 10692 16584
rect 10560 16544 10692 16572
rect 10560 16532 10566 16544
rect 10686 16532 10692 16544
rect 10744 16572 10750 16584
rect 10965 16575 11023 16581
rect 10965 16572 10977 16575
rect 10744 16544 10977 16572
rect 10744 16532 10750 16544
rect 10965 16541 10977 16544
rect 11011 16541 11023 16575
rect 10965 16535 11023 16541
rect 11072 16544 11560 16572
rect 11072 16504 11100 16544
rect 10336 16476 11100 16504
rect 11232 16507 11290 16513
rect 11232 16473 11244 16507
rect 11278 16504 11290 16507
rect 11422 16504 11428 16516
rect 11278 16476 11428 16504
rect 11278 16473 11290 16476
rect 11232 16467 11290 16473
rect 10284 16464 10290 16467
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 11532 16504 11560 16544
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 14274 16572 14280 16584
rect 11756 16544 14280 16572
rect 11756 16532 11762 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15010 16532 15016 16584
rect 15068 16572 15074 16584
rect 15948 16572 15976 16612
rect 16761 16609 16773 16612
rect 16807 16609 16819 16643
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 16761 16603 16819 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 15068 16544 15976 16572
rect 16025 16575 16083 16581
rect 15068 16532 15074 16544
rect 16025 16541 16037 16575
rect 16071 16572 16083 16575
rect 16206 16572 16212 16584
rect 16071 16544 16212 16572
rect 16071 16541 16083 16544
rect 16025 16535 16083 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17126 16572 17132 16584
rect 17083 16544 17132 16572
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 17402 16532 17408 16584
rect 17460 16572 17466 16584
rect 17770 16572 17776 16584
rect 17460 16544 17505 16572
rect 17731 16544 17776 16572
rect 17460 16532 17466 16544
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18322 16572 18328 16584
rect 18283 16544 18328 16572
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 12342 16504 12348 16516
rect 11532 16476 12348 16504
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 13262 16504 13268 16516
rect 13223 16476 13268 16504
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 13906 16464 13912 16516
rect 13964 16504 13970 16516
rect 15286 16504 15292 16516
rect 13964 16476 15292 16504
rect 13964 16464 13970 16476
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 15780 16507 15838 16513
rect 15780 16473 15792 16507
rect 15826 16504 15838 16507
rect 16114 16504 16120 16516
rect 15826 16476 16120 16504
rect 15826 16473 15838 16476
rect 15780 16467 15838 16473
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 7340 16408 7503 16436
rect 7340 16396 7346 16408
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 8294 16436 8300 16448
rect 7708 16408 8300 16436
rect 7708 16396 7714 16408
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 8573 16439 8631 16445
rect 8573 16436 8585 16439
rect 8444 16408 8585 16436
rect 8444 16396 8450 16408
rect 8573 16405 8585 16408
rect 8619 16405 8631 16439
rect 8573 16399 8631 16405
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9582 16436 9588 16448
rect 9171 16408 9588 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11790 16436 11796 16448
rect 11020 16408 11796 16436
rect 11020 16396 11026 16408
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 12802 16436 12808 16448
rect 12763 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 14642 16436 14648 16448
rect 14603 16408 14648 16436
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 3878 16232 3884 16244
rect 3007 16204 3884 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 3878 16192 3884 16204
rect 3936 16232 3942 16244
rect 4522 16232 4528 16244
rect 3936 16204 4528 16232
rect 3936 16192 3942 16204
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 4985 16235 5043 16241
rect 4985 16201 4997 16235
rect 5031 16232 5043 16235
rect 5994 16232 6000 16244
rect 5031 16204 6000 16232
rect 5031 16201 5043 16204
rect 4985 16195 5043 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 6972 16204 10149 16232
rect 6972 16192 6978 16204
rect 10137 16201 10149 16204
rect 10183 16232 10195 16235
rect 10962 16232 10968 16244
rect 10183 16204 10968 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 12621 16235 12679 16241
rect 12621 16232 12633 16235
rect 11204 16204 12633 16232
rect 11204 16192 11210 16204
rect 12621 16201 12633 16204
rect 12667 16201 12679 16235
rect 14550 16232 14556 16244
rect 12621 16195 12679 16201
rect 14200 16204 14556 16232
rect 3326 16124 3332 16176
rect 3384 16164 3390 16176
rect 3384 16136 4108 16164
rect 3384 16124 3390 16136
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1670 16096 1676 16108
rect 1627 16068 1676 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 1848 16099 1906 16105
rect 1848 16065 1860 16099
rect 1894 16096 1906 16099
rect 2222 16096 2228 16108
rect 1894 16068 2228 16096
rect 1894 16065 1906 16068
rect 1848 16059 1906 16065
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 3602 16096 3608 16108
rect 3563 16068 3608 16096
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 3712 16028 3740 16059
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3936 16068 3985 16096
rect 3936 16056 3942 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 4080 16096 4108 16136
rect 4338 16124 4344 16176
rect 4396 16164 4402 16176
rect 4801 16167 4859 16173
rect 4801 16164 4813 16167
rect 4396 16136 4813 16164
rect 4396 16124 4402 16136
rect 4801 16133 4813 16136
rect 4847 16133 4859 16167
rect 4801 16127 4859 16133
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 7101 16167 7159 16173
rect 7101 16164 7113 16167
rect 6604 16136 7113 16164
rect 6604 16124 6610 16136
rect 7101 16133 7113 16136
rect 7147 16164 7159 16167
rect 7282 16164 7288 16176
rect 7147 16136 7288 16164
rect 7147 16133 7159 16136
rect 7101 16127 7159 16133
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 7650 16124 7656 16176
rect 7708 16164 7714 16176
rect 8018 16173 8024 16176
rect 7929 16167 7987 16173
rect 7929 16164 7941 16167
rect 7708 16136 7941 16164
rect 7708 16124 7714 16136
rect 7929 16133 7941 16136
rect 7975 16133 7987 16167
rect 7929 16127 7987 16133
rect 8017 16127 8024 16173
rect 8076 16164 8082 16176
rect 8076 16136 8117 16164
rect 8018 16124 8024 16127
rect 8076 16124 8082 16136
rect 8294 16124 8300 16176
rect 8352 16164 8358 16176
rect 12250 16164 12256 16176
rect 8352 16136 12256 16164
rect 8352 16124 8358 16136
rect 4706 16096 4712 16108
rect 4080 16068 4712 16096
rect 3973 16059 4031 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7765 16099 7823 16105
rect 7765 16096 7777 16099
rect 7248 16068 7777 16096
rect 7248 16056 7254 16068
rect 7765 16065 7777 16068
rect 7811 16065 7823 16099
rect 7765 16059 7823 16065
rect 8159 16099 8217 16105
rect 8159 16065 8171 16099
rect 8205 16096 8217 16099
rect 8205 16068 8340 16096
rect 8205 16065 8217 16068
rect 8159 16059 8217 16065
rect 8312 16040 8340 16068
rect 8662 16056 8668 16108
rect 8720 16096 8726 16108
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 8720 16068 8769 16096
rect 8720 16056 8726 16068
rect 8757 16065 8769 16068
rect 8803 16096 8815 16099
rect 8846 16096 8852 16108
rect 8803 16068 8852 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9030 16105 9036 16108
rect 9024 16059 9036 16105
rect 9088 16096 9094 16108
rect 9088 16068 9124 16096
rect 9030 16056 9036 16059
rect 9088 16056 9094 16068
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 10778 16096 10784 16108
rect 9640 16068 10640 16096
rect 10739 16068 10784 16096
rect 9640 16056 9646 16068
rect 3620 16000 3740 16028
rect 3620 15972 3648 16000
rect 4062 15988 4068 16040
rect 4120 16028 4126 16040
rect 5445 16031 5503 16037
rect 5445 16028 5457 16031
rect 4120 16000 5457 16028
rect 4120 15988 4126 16000
rect 5445 15997 5457 16000
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 5718 15988 5724 16040
rect 5776 16028 5782 16040
rect 5905 16031 5963 16037
rect 5905 16028 5917 16031
rect 5776 16000 5917 16028
rect 5776 15988 5782 16000
rect 5905 15997 5917 16000
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 8294 15988 8300 16040
rect 8352 15988 8358 16040
rect 10612 16028 10640 16068
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 10888 16028 10916 16059
rect 11072 16037 11100 16136
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 12406 16136 12848 16164
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11514 16096 11520 16108
rect 11195 16068 11520 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 12406 16096 12434 16136
rect 12820 16105 12848 16136
rect 13446 16124 13452 16176
rect 13504 16164 13510 16176
rect 14200 16173 14228 16204
rect 14550 16192 14556 16204
rect 14608 16232 14614 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 14608 16204 16313 16232
rect 14608 16192 14614 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 16301 16195 16359 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 13504 16136 14105 16164
rect 13504 16124 13510 16136
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 14093 16127 14151 16133
rect 14185 16167 14243 16173
rect 14185 16133 14197 16167
rect 14231 16133 14243 16167
rect 14185 16127 14243 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 15166 16167 15224 16173
rect 15166 16164 15178 16167
rect 14424 16136 15178 16164
rect 14424 16124 14430 16136
rect 15166 16133 15178 16136
rect 15212 16133 15224 16167
rect 15166 16127 15224 16133
rect 15378 16124 15384 16176
rect 15436 16164 15442 16176
rect 17190 16167 17248 16173
rect 17190 16164 17202 16167
rect 15436 16136 17202 16164
rect 15436 16124 15442 16136
rect 17190 16133 17202 16136
rect 17236 16133 17248 16167
rect 17190 16127 17248 16133
rect 17402 16124 17408 16176
rect 17460 16124 17466 16176
rect 11716 16068 12434 16096
rect 12805 16099 12863 16105
rect 10612 16000 10916 16028
rect 3602 15920 3608 15972
rect 3660 15960 3666 15972
rect 4246 15960 4252 15972
rect 3660 15932 4252 15960
rect 3660 15920 3666 15932
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 4430 15960 4436 15972
rect 4391 15932 4436 15960
rect 4430 15920 4436 15932
rect 4488 15920 4494 15972
rect 4982 15960 4988 15972
rect 4540 15932 4988 15960
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 3421 15895 3479 15901
rect 3421 15892 3433 15895
rect 3108 15864 3433 15892
rect 3108 15852 3114 15864
rect 3421 15861 3433 15864
rect 3467 15861 3479 15895
rect 3421 15855 3479 15861
rect 3694 15852 3700 15904
rect 3752 15892 3758 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 3752 15864 3893 15892
rect 3752 15852 3758 15864
rect 3881 15861 3893 15864
rect 3927 15861 3939 15895
rect 3881 15855 3939 15861
rect 3970 15852 3976 15904
rect 4028 15892 4034 15904
rect 4540 15892 4568 15932
rect 4982 15920 4988 15932
rect 5040 15920 5046 15972
rect 5166 15920 5172 15972
rect 5224 15960 5230 15972
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 5224 15932 5641 15960
rect 5224 15920 5230 15932
rect 5629 15929 5641 15932
rect 5675 15960 5687 15963
rect 6086 15960 6092 15972
rect 5675 15932 6092 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 6733 15963 6791 15969
rect 6733 15929 6745 15963
rect 6779 15960 6791 15963
rect 6822 15960 6828 15972
rect 6779 15932 6828 15960
rect 6779 15929 6791 15932
rect 6733 15923 6791 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 10888 15960 10916 16000
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11716 15960 11744 16068
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11940 16000 12173 16028
rect 11940 15988 11946 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12161 15991 12219 15997
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 12894 16028 12900 16040
rect 12308 16000 12900 16028
rect 12308 15988 12314 16000
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 8402 15932 8800 15960
rect 10888 15932 11744 15960
rect 4798 15892 4804 15904
rect 4028 15864 4568 15892
rect 4759 15864 4804 15892
rect 4028 15852 4034 15864
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7834 15892 7840 15904
rect 7331 15864 7840 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8297 15895 8355 15901
rect 8297 15861 8309 15895
rect 8343 15892 8355 15895
rect 8402 15892 8430 15932
rect 8343 15864 8430 15892
rect 8772 15892 8800 15932
rect 11790 15920 11796 15972
rect 11848 15960 11854 15972
rect 13004 15960 13032 16059
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13909 16099 13967 16105
rect 13136 16068 13229 16096
rect 13136 16056 13142 16068
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 14277 16099 14335 16105
rect 13955 16068 14044 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 11848 15932 13032 15960
rect 11848 15920 11854 15932
rect 9490 15892 9496 15904
rect 8772 15864 9496 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11698 15892 11704 15904
rect 11659 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 13096 15892 13124 16056
rect 13170 15920 13176 15972
rect 13228 15960 13234 15972
rect 14016 15960 14044 16068
rect 14277 16065 14289 16099
rect 14323 16065 14335 16099
rect 16298 16096 16304 16108
rect 14277 16059 14335 16065
rect 14384 16068 16304 16096
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14292 16028 14320 16059
rect 14148 16000 14320 16028
rect 14148 15988 14154 16000
rect 14384 15960 14412 16068
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17420 16096 17448 16124
rect 17052 16068 17448 16096
rect 14918 16028 14924 16040
rect 14879 16000 14924 16028
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 15930 15988 15936 16040
rect 15988 16028 15994 16040
rect 17052 16028 17080 16068
rect 15988 16000 17080 16028
rect 15988 15988 15994 16000
rect 13228 15932 14412 15960
rect 13228 15920 13234 15932
rect 12492 15864 13124 15892
rect 14461 15895 14519 15901
rect 12492 15852 12498 15864
rect 14461 15861 14473 15895
rect 14507 15892 14519 15895
rect 14734 15892 14740 15904
rect 14507 15864 14740 15892
rect 14507 15861 14519 15864
rect 14461 15855 14519 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 16850 15892 16856 15904
rect 14976 15864 16856 15892
rect 14976 15852 14982 15864
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 18046 15852 18052 15904
rect 18104 15892 18110 15904
rect 19242 15892 19248 15904
rect 18104 15864 19248 15892
rect 18104 15852 18110 15864
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 1544 15660 4016 15688
rect 1544 15648 1550 15660
rect 658 15580 664 15632
rect 716 15620 722 15632
rect 716 15592 3832 15620
rect 716 15580 722 15592
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15521 2467 15555
rect 3050 15552 3056 15564
rect 2409 15515 2467 15521
rect 2516 15524 3056 15552
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 2424 15416 2452 15515
rect 2516 15493 2544 15524
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 3694 15552 3700 15564
rect 3436 15524 3700 15552
rect 3436 15493 3464 15524
rect 3694 15512 3700 15524
rect 3752 15512 3758 15564
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3421 15487 3479 15493
rect 3007 15456 3096 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3068 15428 3096 15456
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3804 15484 3832 15592
rect 3988 15561 4016 15660
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 4948 15660 6132 15688
rect 4948 15648 4954 15660
rect 3973 15555 4031 15561
rect 3973 15521 3985 15555
rect 4019 15521 4031 15555
rect 3973 15515 4031 15521
rect 4229 15487 4287 15493
rect 4229 15484 4241 15487
rect 3804 15456 4241 15484
rect 3421 15447 3479 15453
rect 4229 15453 4241 15456
rect 4275 15453 4287 15487
rect 4229 15447 4287 15453
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 6104 15493 6132 15660
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 7558 15688 7564 15700
rect 7156 15660 7564 15688
rect 7156 15648 7162 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 9122 15688 9128 15700
rect 7944 15660 9128 15688
rect 7282 15580 7288 15632
rect 7340 15620 7346 15632
rect 7377 15623 7435 15629
rect 7377 15620 7389 15623
rect 7340 15592 7389 15620
rect 7340 15580 7346 15592
rect 7377 15589 7389 15592
rect 7423 15620 7435 15623
rect 7834 15620 7840 15632
rect 7423 15592 7840 15620
rect 7423 15589 7435 15592
rect 7377 15583 7435 15589
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 7944 15552 7972 15660
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 11241 15691 11299 15697
rect 9272 15660 10548 15688
rect 9272 15648 9278 15660
rect 10520 15632 10548 15660
rect 11241 15657 11253 15691
rect 11287 15657 11299 15691
rect 11241 15651 11299 15657
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 8076 15592 8340 15620
rect 8076 15580 8082 15592
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 6512 15524 8125 15552
rect 6512 15512 6518 15524
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 8312 15552 8340 15592
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 8754 15620 8760 15632
rect 8444 15592 8760 15620
rect 8444 15580 8450 15592
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 10502 15580 10508 15632
rect 10560 15580 10566 15632
rect 11256 15620 11284 15651
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12768 15660 12909 15688
rect 12768 15648 12774 15660
rect 12897 15657 12909 15660
rect 12943 15657 12955 15691
rect 12897 15651 12955 15657
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 13320 15660 14289 15688
rect 13320 15648 13326 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15010 15688 15016 15700
rect 14884 15660 15016 15688
rect 14884 15648 14890 15660
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15378 15688 15384 15700
rect 15120 15660 15384 15688
rect 11072 15592 11284 15620
rect 11885 15623 11943 15629
rect 8938 15552 8944 15564
rect 8312 15524 8944 15552
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5132 15456 5825 15484
rect 5132 15444 5138 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6788 15456 7696 15484
rect 6788 15444 6794 15456
rect 2424 15388 2728 15416
rect 1857 15351 1915 15357
rect 1857 15317 1869 15351
rect 1903 15348 1915 15351
rect 1946 15348 1952 15360
rect 1903 15320 1952 15348
rect 1903 15317 1915 15320
rect 1857 15311 1915 15317
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 2700 15348 2728 15388
rect 3050 15376 3056 15428
rect 3108 15416 3114 15428
rect 3878 15416 3884 15428
rect 3108 15388 3884 15416
rect 3108 15376 3114 15388
rect 3878 15376 3884 15388
rect 3936 15376 3942 15428
rect 6273 15419 6331 15425
rect 6273 15416 6285 15419
rect 4356 15388 6285 15416
rect 4356 15348 4384 15388
rect 6273 15385 6285 15388
rect 6319 15385 6331 15419
rect 6273 15379 6331 15385
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 7101 15419 7159 15425
rect 7101 15416 7113 15419
rect 6972 15388 7113 15416
rect 6972 15376 6978 15388
rect 7101 15385 7113 15388
rect 7147 15385 7159 15419
rect 7668 15416 7696 15456
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 8312 15493 8340 15524
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 11072 15552 11100 15592
rect 11885 15589 11897 15623
rect 11931 15620 11943 15623
rect 12158 15620 12164 15632
rect 11931 15592 12164 15620
rect 11931 15589 11943 15592
rect 11885 15583 11943 15589
rect 12158 15580 12164 15592
rect 12216 15580 12222 15632
rect 13538 15620 13544 15632
rect 13499 15592 13544 15620
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 15120 15620 15148 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 15473 15691 15531 15697
rect 15473 15657 15485 15691
rect 15519 15688 15531 15691
rect 15930 15688 15936 15700
rect 15519 15660 15936 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16301 15691 16359 15697
rect 16301 15657 16313 15691
rect 16347 15688 16359 15691
rect 17862 15688 17868 15700
rect 16347 15660 17868 15688
rect 16347 15657 16359 15660
rect 16301 15651 16359 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 15286 15620 15292 15632
rect 14056 15592 15148 15620
rect 15203 15592 15292 15620
rect 14056 15580 14062 15592
rect 10428 15524 11100 15552
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7800 15456 8033 15484
rect 7800 15444 7806 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8296 15487 8354 15493
rect 8296 15453 8308 15487
rect 8342 15453 8354 15487
rect 8296 15447 8354 15453
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 9674 15484 9680 15496
rect 8619 15456 9680 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 8110 15416 8116 15428
rect 7668 15388 8116 15416
rect 7101 15379 7159 15385
rect 8110 15376 8116 15388
rect 8168 15416 8174 15428
rect 8404 15416 8432 15447
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10428 15484 10456 15524
rect 10152 15456 10456 15484
rect 10505 15487 10563 15493
rect 8168 15388 8432 15416
rect 8168 15376 8174 15388
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 10152 15416 10180 15456
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 10686 15484 10692 15496
rect 10551 15456 10692 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 8812 15388 10180 15416
rect 10260 15419 10318 15425
rect 8812 15376 8818 15388
rect 10260 15385 10272 15419
rect 10306 15416 10318 15419
rect 10870 15416 10876 15428
rect 10306 15388 10876 15416
rect 10306 15385 10318 15388
rect 10260 15379 10318 15385
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 2700 15320 4384 15348
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 5353 15351 5411 15357
rect 5353 15348 5365 15351
rect 5224 15320 5365 15348
rect 5224 15308 5230 15320
rect 5353 15317 5365 15320
rect 5399 15317 5411 15351
rect 5353 15311 5411 15317
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 5905 15351 5963 15357
rect 5905 15348 5917 15351
rect 5868 15320 5917 15348
rect 5868 15308 5874 15320
rect 5905 15317 5917 15320
rect 5951 15317 5963 15351
rect 5905 15311 5963 15317
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 7190 15348 7196 15360
rect 6696 15320 7196 15348
rect 6696 15308 6702 15320
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 7561 15351 7619 15357
rect 7561 15317 7573 15351
rect 7607 15348 7619 15351
rect 8938 15348 8944 15360
rect 7607 15320 8944 15348
rect 7607 15317 7619 15320
rect 7561 15311 7619 15317
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15348 9370 15360
rect 10686 15348 10692 15360
rect 9364 15320 10692 15348
rect 9364 15308 9370 15320
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11072 15348 11100 15524
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 12066 15552 12072 15564
rect 11296 15524 12072 15552
rect 11296 15512 11302 15524
rect 12066 15512 12072 15524
rect 12124 15552 12130 15564
rect 12710 15552 12716 15564
rect 12124 15524 12716 15552
rect 12124 15512 12130 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13044 15524 14504 15552
rect 13044 15512 13050 15524
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 13262 15484 13268 15496
rect 11471 15480 12572 15484
rect 12636 15480 13268 15484
rect 11471 15456 13268 15480
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 12544 15452 12664 15456
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 11790 15376 11796 15428
rect 11848 15416 11854 15428
rect 12069 15419 12127 15425
rect 12069 15416 12081 15419
rect 11848 15388 12081 15416
rect 11848 15376 11854 15388
rect 12069 15385 12081 15388
rect 12115 15385 12127 15419
rect 12069 15379 12127 15385
rect 12253 15419 12311 15425
rect 12253 15385 12265 15419
rect 12299 15416 12311 15419
rect 12434 15416 12440 15428
rect 12299 15388 12440 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 12268 15348 12296 15379
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 12865 15419 12923 15425
rect 12865 15416 12877 15419
rect 12544 15388 12877 15416
rect 12544 15360 12572 15388
rect 12865 15385 12877 15388
rect 12911 15385 12923 15419
rect 12865 15379 12923 15385
rect 12986 15376 12992 15428
rect 13044 15416 13050 15428
rect 13081 15419 13139 15425
rect 13081 15416 13093 15419
rect 13044 15388 13093 15416
rect 13044 15376 13050 15388
rect 13081 15385 13093 15388
rect 13127 15385 13139 15419
rect 13081 15379 13139 15385
rect 13648 15360 13676 15524
rect 14476 15493 14504 15524
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 15203 15552 15231 15592
rect 15286 15580 15292 15592
rect 15344 15580 15350 15632
rect 18046 15580 18052 15632
rect 18104 15620 18110 15632
rect 18325 15623 18383 15629
rect 18325 15620 18337 15623
rect 18104 15592 18337 15620
rect 18104 15580 18110 15592
rect 18325 15589 18337 15592
rect 18371 15589 18383 15623
rect 18325 15583 18383 15589
rect 14608 15524 15231 15552
rect 14608 15512 14614 15524
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15486 14979 15487
rect 15010 15486 15016 15496
rect 14967 15458 15016 15486
rect 14967 15453 14979 15458
rect 14921 15447 14979 15453
rect 15010 15444 15016 15458
rect 15068 15444 15074 15496
rect 15203 15493 15231 15524
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15930 15484 15936 15496
rect 15891 15456 15936 15484
rect 15289 15447 15347 15453
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15302 15416 15330 15447
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16942 15484 16948 15496
rect 16264 15456 16948 15484
rect 16264 15444 16270 15456
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17770 15484 17776 15496
rect 17144 15456 17776 15484
rect 14148 15388 15330 15416
rect 16301 15419 16359 15425
rect 14148 15376 14154 15388
rect 16301 15385 16313 15419
rect 16347 15416 16359 15419
rect 16850 15416 16856 15428
rect 16347 15388 16856 15416
rect 16347 15385 16359 15388
rect 16301 15379 16359 15385
rect 16850 15376 16856 15388
rect 16908 15416 16914 15428
rect 17144 15416 17172 15456
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 17218 15425 17224 15428
rect 16908 15388 17172 15416
rect 16908 15376 16914 15388
rect 17212 15379 17224 15425
rect 17276 15416 17282 15428
rect 18414 15416 18420 15428
rect 17276 15388 17312 15416
rect 18248 15388 18420 15416
rect 17218 15376 17224 15379
rect 17276 15376 17282 15388
rect 11072 15320 12296 15348
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 12710 15348 12716 15360
rect 12671 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 13630 15308 13636 15360
rect 13688 15308 13694 15360
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 15746 15348 15752 15360
rect 13780 15320 15752 15348
rect 13780 15308 13786 15320
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 18248 15348 18276 15388
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 16531 15320 18276 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3602 15144 3608 15156
rect 3007 15116 3608 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3602 15104 3608 15116
rect 3660 15144 3666 15156
rect 4890 15144 4896 15156
rect 3660 15116 4896 15144
rect 3660 15104 3666 15116
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 5074 15144 5080 15156
rect 5035 15116 5080 15144
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 8754 15144 8760 15156
rect 5184 15116 8760 15144
rect 3615 15048 4936 15076
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 1670 15008 1676 15020
rect 1627 14980 1676 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 1848 15011 1906 15017
rect 1848 14977 1860 15011
rect 1894 15008 1906 15011
rect 2314 15008 2320 15020
rect 1894 14980 2320 15008
rect 1894 14977 1906 14980
rect 1848 14971 1906 14977
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 3615 15017 3643 15048
rect 3600 15011 3658 15017
rect 3600 14977 3612 15011
rect 3646 14977 3658 15011
rect 3600 14971 3658 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 3712 14940 3740 14971
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 3970 15008 3976 15020
rect 3844 14980 3889 15008
rect 3931 14980 3976 15008
rect 3844 14968 3850 14980
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4522 15008 4528 15020
rect 4120 14980 4165 15008
rect 4483 14980 4528 15008
rect 4120 14968 4126 14980
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 4908 15017 4936 15048
rect 4982 15036 4988 15088
rect 5040 15076 5046 15088
rect 5184 15076 5212 15116
rect 5534 15076 5540 15088
rect 5040 15048 5212 15076
rect 5495 15048 5540 15076
rect 5040 15036 5046 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 5753 15079 5811 15085
rect 5753 15045 5765 15079
rect 5799 15076 5811 15079
rect 5994 15076 6000 15088
rect 5799 15048 6000 15076
rect 5799 15045 5811 15048
rect 5753 15039 5811 15045
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 6840 15085 6868 15116
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9769 15147 9827 15153
rect 9769 15144 9781 15147
rect 9456 15116 9781 15144
rect 9456 15104 9462 15116
rect 9769 15113 9781 15116
rect 9815 15113 9827 15147
rect 10778 15144 10784 15156
rect 9769 15107 9827 15113
rect 9968 15116 10784 15144
rect 6825 15079 6883 15085
rect 6825 15045 6837 15079
rect 6871 15045 6883 15079
rect 6825 15039 6883 15045
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 7805 15079 7863 15085
rect 7805 15076 7817 15079
rect 7340 15048 7817 15076
rect 7340 15036 7346 15048
rect 7805 15045 7817 15048
rect 7851 15045 7863 15079
rect 7805 15039 7863 15045
rect 8021 15079 8079 15085
rect 8021 15045 8033 15079
rect 8067 15076 8079 15079
rect 8110 15076 8116 15088
rect 8067 15048 8116 15076
rect 8067 15045 8079 15048
rect 8021 15039 8079 15045
rect 8110 15036 8116 15048
rect 8168 15036 8174 15088
rect 8294 15036 8300 15088
rect 8352 15076 8358 15088
rect 9858 15076 9864 15088
rect 8352 15048 9864 15076
rect 8352 15036 8358 15048
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5350 15008 5356 15020
rect 4939 14980 5356 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 4816 14940 4844 14971
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 9674 15008 9680 15020
rect 8895 14980 9680 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 5074 14940 5080 14952
rect 3712 14912 5080 14940
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 7024 14940 7052 14971
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9968 15017 9996 15116
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 12802 15144 12808 15156
rect 11072 15116 12808 15144
rect 10137 15079 10195 15085
rect 10137 15045 10149 15079
rect 10183 15076 10195 15079
rect 10962 15076 10968 15088
rect 10183 15048 10968 15076
rect 10183 15045 10195 15048
rect 10137 15039 10195 15045
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 9948 15011 10006 15017
rect 9948 14977 9960 15011
rect 9994 14977 10006 15011
rect 9948 14971 10006 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10320 15011 10378 15017
rect 10320 14977 10332 15011
rect 10366 14977 10378 15011
rect 10320 14971 10378 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 11072 15008 11100 15116
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 15930 15144 15936 15156
rect 14608 15116 15936 15144
rect 14608 15104 14614 15116
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 17402 15104 17408 15156
rect 17460 15144 17466 15156
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 17460 15116 18337 15144
rect 17460 15104 17466 15116
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 11869 15079 11927 15085
rect 11869 15045 11881 15079
rect 11915 15076 11927 15079
rect 12066 15076 12072 15088
rect 11915 15045 11928 15076
rect 12027 15048 12072 15076
rect 11869 15039 11928 15045
rect 10459 14980 11100 15008
rect 11149 15011 11207 15017
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11238 15008 11244 15020
rect 11195 14980 11244 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 8018 14940 8024 14952
rect 5500 14912 5948 14940
rect 7024 14912 8024 14940
rect 5500 14900 5506 14912
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14872 3479 14875
rect 5810 14872 5816 14884
rect 3467 14844 5816 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 5810 14832 5816 14844
rect 5868 14832 5874 14884
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 5920 14813 5948 14912
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8168 14912 8769 14940
rect 8168 14900 8174 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 10060 14940 10088 14971
rect 9640 14912 10088 14940
rect 10336 14940 10364 14971
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 11698 14940 11704 14952
rect 10336 14912 11704 14940
rect 9640 14900 9646 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7558 14872 7564 14884
rect 7239 14844 7564 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 10502 14872 10508 14884
rect 8036 14844 10508 14872
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 4948 14776 5733 14804
rect 4948 14764 4954 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6730 14804 6736 14816
rect 5951 14776 6736 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7653 14807 7711 14813
rect 7653 14804 7665 14807
rect 7524 14776 7665 14804
rect 7524 14764 7530 14776
rect 7653 14773 7665 14776
rect 7699 14773 7711 14807
rect 7653 14767 7711 14773
rect 7837 14807 7895 14813
rect 7837 14773 7849 14807
rect 7883 14804 7895 14807
rect 8036 14804 8064 14844
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 10686 14832 10692 14884
rect 10744 14872 10750 14884
rect 11900 14872 11928 15039
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 13170 15036 13176 15088
rect 13228 15076 13234 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13228 15048 13369 15076
rect 13228 15036 13234 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 14169 15079 14227 15085
rect 14169 15045 14181 15079
rect 14215 15045 14227 15079
rect 14169 15039 14227 15045
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 12032 14980 12541 15008
rect 12032 14968 12038 14980
rect 12529 14977 12541 14980
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 14184 15008 14212 15039
rect 14340 15036 14346 15088
rect 14398 15076 14404 15088
rect 16298 15076 16304 15088
rect 14398 15048 14443 15076
rect 15764 15048 16304 15076
rect 14398 15036 14404 15048
rect 15764 15020 15792 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 17190 15079 17248 15085
rect 17190 15045 17202 15079
rect 17236 15076 17248 15079
rect 17770 15076 17776 15088
rect 17236 15048 17776 15076
rect 17236 15045 17248 15048
rect 17190 15039 17248 15045
rect 17770 15036 17776 15048
rect 17828 15036 17834 15088
rect 13587 14980 14044 15008
rect 14184 14980 15700 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 14016 14881 14044 14980
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15562 14940 15568 14952
rect 14875 14912 15568 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 15672 14940 15700 14980
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16025 15011 16083 15017
rect 15804 14980 15897 15008
rect 15804 14968 15810 14980
rect 16025 14977 16037 15011
rect 16071 14977 16083 15011
rect 16025 14971 16083 14977
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16206 15008 16212 15020
rect 16163 14980 16212 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16040 14940 16068 14971
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 18046 15008 18052 15020
rect 16868 14980 18052 15008
rect 16868 14940 16896 14980
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 15672 14912 16896 14940
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 17000 14912 17045 14940
rect 17000 14900 17006 14912
rect 10744 14844 11928 14872
rect 14001 14875 14059 14881
rect 10744 14832 10750 14844
rect 14001 14841 14013 14875
rect 14047 14872 14059 14875
rect 14550 14872 14556 14884
rect 14047 14844 14556 14872
rect 14047 14841 14059 14844
rect 14001 14835 14059 14841
rect 14550 14832 14556 14844
rect 14608 14832 14614 14884
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14841 15255 14875
rect 15197 14835 15255 14841
rect 15289 14875 15347 14881
rect 15289 14841 15301 14875
rect 15335 14872 15347 14875
rect 15335 14844 16988 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 8570 14804 8576 14816
rect 7883 14776 8064 14804
rect 8531 14776 8576 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 8904 14776 10977 14804
rect 8904 14764 8910 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 10965 14767 11023 14773
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 11204 14776 11713 14804
rect 11204 14764 11210 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11848 14776 11897 14804
rect 11848 14764 11854 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 11885 14767 11943 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 14185 14807 14243 14813
rect 14185 14773 14197 14807
rect 14231 14804 14243 14807
rect 14642 14804 14648 14816
rect 14231 14776 14648 14804
rect 14231 14773 14243 14776
rect 14185 14767 14243 14773
rect 14642 14764 14648 14776
rect 14700 14804 14706 14816
rect 15212 14804 15240 14835
rect 15378 14804 15384 14816
rect 14700 14776 15384 14804
rect 14700 14764 14706 14776
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 15838 14804 15844 14816
rect 15799 14776 15844 14804
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 16301 14807 16359 14813
rect 16301 14773 16313 14807
rect 16347 14804 16359 14807
rect 16390 14804 16396 14816
rect 16347 14776 16396 14804
rect 16347 14773 16359 14776
rect 16301 14767 16359 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16960 14804 16988 14844
rect 18138 14804 18144 14816
rect 16960 14776 18144 14804
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 750 14560 756 14612
rect 808 14600 814 14612
rect 808 14572 2544 14600
rect 808 14560 814 14572
rect 2516 14532 2544 14572
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3936 14572 4169 14600
rect 3936 14560 3942 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 4430 14560 4436 14612
rect 4488 14600 4494 14612
rect 5166 14600 5172 14612
rect 4488 14572 5172 14600
rect 4488 14560 4494 14572
rect 5166 14560 5172 14572
rect 5224 14600 5230 14612
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 5224 14572 5825 14600
rect 5224 14560 5230 14572
rect 5813 14569 5825 14572
rect 5859 14569 5871 14603
rect 5813 14563 5871 14569
rect 6825 14603 6883 14609
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7282 14600 7288 14612
rect 6871 14572 7288 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 8386 14600 8392 14612
rect 7392 14572 8392 14600
rect 3973 14535 4031 14541
rect 3973 14532 3985 14535
rect 2516 14504 3985 14532
rect 3973 14501 3985 14504
rect 4019 14501 4031 14535
rect 3973 14495 4031 14501
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 5442 14532 5448 14544
rect 4672 14504 5448 14532
rect 4672 14492 4678 14504
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 5902 14492 5908 14544
rect 5960 14532 5966 14544
rect 7392 14532 7420 14572
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 9309 14603 9367 14609
rect 9309 14569 9321 14603
rect 9355 14600 9367 14603
rect 10318 14600 10324 14612
rect 9355 14572 10324 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 11238 14600 11244 14612
rect 10560 14572 11244 14600
rect 10560 14560 10566 14572
rect 11238 14560 11244 14572
rect 11296 14600 11302 14612
rect 12434 14600 12440 14612
rect 11296 14572 12020 14600
rect 12395 14572 12440 14600
rect 11296 14560 11302 14572
rect 7558 14532 7564 14544
rect 5960 14504 6592 14532
rect 5960 14492 5966 14504
rect 4982 14464 4988 14476
rect 2746 14436 4988 14464
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 1670 14396 1676 14408
rect 1627 14368 1676 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 1848 14331 1906 14337
rect 1848 14297 1860 14331
rect 1894 14328 1906 14331
rect 2746 14328 2774 14436
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5534 14424 5540 14476
rect 5592 14464 5598 14476
rect 6181 14467 6239 14473
rect 6181 14464 6193 14467
rect 5592 14436 6193 14464
rect 5592 14424 5598 14436
rect 6181 14433 6193 14436
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4396 14368 4537 14396
rect 4396 14356 4402 14368
rect 4525 14365 4537 14368
rect 4571 14396 4583 14399
rect 5994 14396 6000 14408
rect 4571 14368 6000 14396
rect 4571 14365 4583 14368
rect 4525 14359 4583 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 1894 14300 2774 14328
rect 1894 14297 1906 14300
rect 1848 14291 1906 14297
rect 3418 14288 3424 14340
rect 3476 14328 3482 14340
rect 5169 14331 5227 14337
rect 3476 14300 5120 14328
rect 3476 14288 3482 14300
rect 2961 14263 3019 14269
rect 2961 14229 2973 14263
rect 3007 14260 3019 14263
rect 3050 14260 3056 14272
rect 3007 14232 3056 14260
rect 3007 14229 3019 14232
rect 2961 14223 3019 14229
rect 3050 14220 3056 14232
rect 3108 14260 3114 14272
rect 3970 14260 3976 14272
rect 3108 14232 3976 14260
rect 3108 14220 3114 14232
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 4985 14263 5043 14269
rect 4985 14260 4997 14263
rect 4580 14232 4997 14260
rect 4580 14220 4586 14232
rect 4985 14229 4997 14232
rect 5031 14229 5043 14263
rect 5092 14260 5120 14300
rect 5169 14297 5181 14331
rect 5215 14328 5227 14331
rect 5258 14328 5264 14340
rect 5215 14300 5264 14328
rect 5215 14297 5227 14300
rect 5169 14291 5227 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 5353 14331 5411 14337
rect 5353 14297 5365 14331
rect 5399 14328 5411 14331
rect 5442 14328 5448 14340
rect 5399 14300 5448 14328
rect 5399 14297 5411 14300
rect 5353 14291 5411 14297
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 5810 14260 5816 14272
rect 5092 14232 5816 14260
rect 4985 14223 5043 14229
rect 5810 14220 5816 14232
rect 5868 14260 5874 14272
rect 6086 14260 6092 14272
rect 5868 14232 6092 14260
rect 5868 14220 5874 14232
rect 6086 14220 6092 14232
rect 6144 14220 6150 14272
rect 6564 14260 6592 14504
rect 6672 14504 7420 14532
rect 7484 14504 7564 14532
rect 6672 14396 6700 14504
rect 6756 14399 6814 14405
rect 6756 14396 6768 14399
rect 6672 14368 6768 14396
rect 6756 14365 6768 14368
rect 6802 14365 6814 14399
rect 6914 14396 6920 14408
rect 6875 14368 6920 14396
rect 6756 14359 6814 14365
rect 6914 14356 6920 14368
rect 6972 14396 6978 14408
rect 7484 14396 7512 14504
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 11992 14532 12020 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13872 14572 14289 14600
rect 13872 14560 13878 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 15010 14560 15016 14612
rect 15068 14600 15074 14612
rect 15194 14600 15200 14612
rect 15068 14572 15200 14600
rect 15068 14560 15074 14572
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 15378 14560 15384 14612
rect 15436 14600 15442 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 15436 14572 15853 14600
rect 15436 14560 15442 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 13078 14532 13084 14544
rect 11992 14504 13084 14532
rect 8202 14464 8208 14476
rect 7576 14436 8208 14464
rect 7576 14405 7604 14436
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 10318 14464 10324 14476
rect 9916 14436 10324 14464
rect 9916 14424 9922 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 11992 14473 12020 14504
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 13170 14492 13176 14544
rect 13228 14532 13234 14544
rect 16868 14532 16896 14563
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17494 14600 17500 14612
rect 17000 14572 17500 14600
rect 17000 14560 17006 14572
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 13228 14504 16896 14532
rect 13228 14492 13234 14504
rect 17126 14492 17132 14544
rect 17184 14532 17190 14544
rect 17221 14535 17279 14541
rect 17221 14532 17233 14535
rect 17184 14504 17233 14532
rect 17184 14492 17190 14504
rect 17221 14501 17233 14504
rect 17267 14501 17279 14535
rect 17221 14495 17279 14501
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 15838 14464 15844 14476
rect 13504 14436 15844 14464
rect 13504 14424 13510 14436
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 16209 14467 16267 14473
rect 15948 14436 16160 14464
rect 6972 14368 7512 14396
rect 7561 14399 7619 14405
rect 6972 14356 6978 14368
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9122 14396 9128 14408
rect 8904 14368 9128 14396
rect 8904 14356 8910 14368
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9490 14396 9496 14408
rect 9451 14368 9496 14396
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 10594 14396 10600 14408
rect 9815 14368 10600 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 13078 14396 13084 14408
rect 13039 14368 13084 14396
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15378 14396 15384 14408
rect 14967 14368 15384 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15620 14368 15761 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 7745 14331 7803 14337
rect 7745 14328 7757 14331
rect 7248 14300 7757 14328
rect 7248 14288 7254 14300
rect 7745 14297 7757 14300
rect 7791 14297 7803 14331
rect 7745 14291 7803 14297
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 6564 14232 7389 14260
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 7760 14260 7788 14291
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8205 14331 8263 14337
rect 8205 14328 8217 14331
rect 7892 14300 8217 14328
rect 7892 14288 7898 14300
rect 8205 14297 8217 14300
rect 8251 14297 8263 14331
rect 8205 14291 8263 14297
rect 8421 14331 8479 14337
rect 8421 14297 8433 14331
rect 8467 14328 8479 14331
rect 9582 14328 9588 14340
rect 8467 14300 9588 14328
rect 8467 14297 8479 14300
rect 8421 14291 8479 14297
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 11698 14328 11704 14340
rect 11756 14337 11762 14340
rect 11668 14300 11704 14328
rect 11698 14288 11704 14300
rect 11756 14291 11768 14337
rect 11756 14288 11762 14291
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 12952 14300 13185 14328
rect 12952 14288 12958 14300
rect 13173 14297 13185 14300
rect 13219 14297 13231 14331
rect 13173 14291 13231 14297
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 15105 14331 15163 14337
rect 15105 14328 15117 14331
rect 14424 14300 15117 14328
rect 14424 14288 14430 14300
rect 15105 14297 15117 14300
rect 15151 14328 15163 14331
rect 15194 14328 15200 14340
rect 15151 14300 15200 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15289 14331 15347 14337
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 15948 14328 15976 14436
rect 15335 14300 15976 14328
rect 16132 14328 16160 14436
rect 16209 14433 16221 14467
rect 16255 14464 16267 14467
rect 16255 14436 18092 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 18064 14405 18092 14436
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 18196 14436 18368 14464
rect 18196 14424 18202 14436
rect 17819 14399 17877 14405
rect 17819 14396 17831 14399
rect 16356 14368 17831 14396
rect 16356 14356 16362 14368
rect 17819 14365 17831 14368
rect 17865 14365 17877 14399
rect 17819 14359 17877 14365
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18230 14396 18236 14408
rect 18191 14368 18236 14396
rect 18049 14359 18107 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18340 14405 18368 14436
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 17957 14331 18015 14337
rect 16132 14300 17908 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 7760 14232 8585 14260
rect 7377 14223 7435 14229
rect 8573 14229 8585 14232
rect 8619 14260 8631 14263
rect 8846 14260 8852 14272
rect 8619 14232 8852 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 9677 14263 9735 14269
rect 9677 14260 9689 14263
rect 9456 14232 9689 14260
rect 9456 14220 9462 14232
rect 9677 14229 9689 14232
rect 9723 14229 9735 14263
rect 9677 14223 9735 14229
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 11238 14260 11244 14272
rect 10643 14232 11244 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 12526 14260 12532 14272
rect 11388 14232 12532 14260
rect 11388 14220 11394 14232
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16264 14232 16681 14260
rect 16264 14220 16270 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16816 14232 16865 14260
rect 16816 14220 16822 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17681 14263 17739 14269
rect 17681 14260 17693 14263
rect 17092 14232 17693 14260
rect 17092 14220 17098 14232
rect 17681 14229 17693 14232
rect 17727 14229 17739 14263
rect 17880 14260 17908 14300
rect 17957 14297 17969 14331
rect 18003 14328 18015 14331
rect 18138 14328 18144 14340
rect 18003 14300 18144 14328
rect 18003 14297 18015 14300
rect 17957 14291 18015 14297
rect 18138 14288 18144 14300
rect 18196 14288 18202 14340
rect 18046 14260 18052 14272
rect 17880 14232 18052 14260
rect 17681 14223 17739 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 18156 14260 18184 14288
rect 18322 14260 18328 14272
rect 18156 14232 18328 14260
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3418 14056 3424 14068
rect 3007 14028 3424 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3878 14056 3884 14068
rect 3839 14028 3884 14056
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 7834 14056 7840 14068
rect 4755 14028 7840 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 9122 14056 9128 14068
rect 8496 14028 9128 14056
rect 8496 14000 8524 14028
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9732 14028 9873 14056
rect 9732 14016 9738 14028
rect 9861 14025 9873 14028
rect 9907 14056 9919 14059
rect 9950 14056 9956 14068
rect 9907 14028 9956 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10321 14059 10379 14065
rect 10321 14056 10333 14059
rect 10192 14028 10333 14056
rect 10192 14016 10198 14028
rect 10321 14025 10333 14028
rect 10367 14056 10379 14059
rect 11330 14056 11336 14068
rect 10367 14028 11336 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11698 14056 11704 14068
rect 11659 14028 11704 14056
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14274 14056 14280 14068
rect 13964 14028 14280 14056
rect 13964 14016 13970 14028
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 14700 14028 15945 14056
rect 14700 14016 14706 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 16632 14028 17785 14056
rect 16632 14016 16638 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 18138 14056 18144 14068
rect 17773 14019 17831 14025
rect 17880 14028 18144 14056
rect 1946 13948 1952 14000
rect 2004 13988 2010 14000
rect 4154 13988 4160 14000
rect 2004 13960 4160 13988
rect 2004 13948 2010 13960
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 4341 13991 4399 13997
rect 4341 13988 4353 13991
rect 4212 13960 4353 13988
rect 4212 13948 4218 13960
rect 4341 13957 4353 13960
rect 4387 13957 4399 13991
rect 4341 13951 4399 13957
rect 4557 13991 4615 13997
rect 4557 13957 4569 13991
rect 4603 13988 4615 13991
rect 5258 13988 5264 14000
rect 4603 13960 5264 13988
rect 4603 13957 4615 13960
rect 4557 13951 4615 13957
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 6794 13991 6852 13997
rect 6794 13988 6806 13991
rect 6288 13960 6806 13988
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 1848 13923 1906 13929
rect 1848 13889 1860 13923
rect 1894 13920 1906 13923
rect 3418 13920 3424 13932
rect 1894 13892 3280 13920
rect 3379 13892 3424 13920
rect 1894 13889 1906 13892
rect 1848 13883 1906 13889
rect 3252 13852 3280 13892
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3697 13923 3755 13929
rect 3568 13892 3613 13920
rect 3568 13880 3574 13892
rect 3697 13889 3709 13923
rect 3743 13920 3755 13923
rect 5074 13920 5080 13932
rect 3743 13892 5080 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 5074 13880 5080 13892
rect 5132 13920 5138 13932
rect 5350 13920 5356 13932
rect 5132 13892 5356 13920
rect 5132 13880 5138 13892
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5523 13923 5581 13929
rect 5523 13889 5535 13923
rect 5569 13920 5581 13923
rect 5569 13892 5764 13920
rect 5569 13889 5581 13892
rect 5523 13883 5581 13889
rect 3252 13824 4109 13852
rect 2590 13744 2596 13796
rect 2648 13784 2654 13796
rect 3786 13784 3792 13796
rect 2648 13756 3792 13784
rect 2648 13744 2654 13756
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 4081 13784 4109 13824
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 5445 13855 5503 13861
rect 5445 13852 5457 13855
rect 4212 13824 5457 13852
rect 4212 13812 4218 13824
rect 5445 13821 5457 13824
rect 5491 13852 5503 13855
rect 5626 13852 5632 13864
rect 5491 13824 5632 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 5074 13784 5080 13796
rect 4081 13756 5080 13784
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 4522 13716 4528 13728
rect 4483 13688 4528 13716
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 5736 13716 5764 13892
rect 5813 13787 5871 13793
rect 5813 13753 5825 13787
rect 5859 13784 5871 13787
rect 6288 13784 6316 13960
rect 6794 13957 6806 13960
rect 6840 13957 6852 13991
rect 6794 13951 6852 13957
rect 6914 13948 6920 14000
rect 6972 13948 6978 14000
rect 8478 13948 8484 14000
rect 8536 13948 8542 14000
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 8726 13991 8784 13997
rect 8726 13988 8738 13991
rect 8628 13960 8738 13988
rect 8628 13948 8634 13960
rect 8726 13957 8738 13960
rect 8772 13957 8784 13991
rect 8726 13951 8784 13957
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 10473 13991 10531 13997
rect 10473 13988 10485 13991
rect 8904 13960 10485 13988
rect 8904 13948 8910 13960
rect 10473 13957 10485 13960
rect 10519 13957 10531 13991
rect 10473 13951 10531 13957
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 11514 13988 11520 14000
rect 10735 13960 11520 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 6932 13920 6960 13948
rect 6696 13892 6960 13920
rect 6696 13880 6702 13892
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 9122 13920 9128 13932
rect 8260 13892 9128 13920
rect 8260 13880 8266 13892
rect 9122 13880 9128 13892
rect 9180 13920 9186 13932
rect 10704 13920 10732 13951
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 15105 13991 15163 13997
rect 15105 13957 15117 13991
rect 15151 13988 15163 13991
rect 15194 13988 15200 14000
rect 15151 13960 15200 13988
rect 15151 13957 15163 13960
rect 15105 13951 15163 13957
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15321 13991 15379 13997
rect 15321 13957 15333 13991
rect 15367 13988 15379 13991
rect 16101 13991 16159 13997
rect 15367 13960 15516 13988
rect 15367 13957 15379 13960
rect 15321 13951 15379 13957
rect 9180 13892 10732 13920
rect 9180 13880 9186 13892
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11296 13892 12081 13920
rect 11296 13880 11302 13892
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13722 13920 13728 13932
rect 13403 13892 13728 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14182 13880 14188 13932
rect 14240 13920 14246 13932
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 14240 13892 14473 13920
rect 14240 13880 14246 13892
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 15488 13920 15516 13960
rect 16101 13957 16113 13991
rect 16147 13988 16159 13991
rect 16206 13988 16212 14000
rect 16147 13960 16212 13988
rect 16147 13957 16159 13960
rect 16101 13951 16159 13957
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16301 13991 16359 13997
rect 16301 13957 16313 13991
rect 16347 13988 16359 13991
rect 16482 13988 16488 14000
rect 16347 13960 16488 13988
rect 16347 13957 16359 13960
rect 16301 13951 16359 13957
rect 16482 13948 16488 13960
rect 16540 13948 16546 14000
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 17000 13960 17325 13988
rect 17000 13948 17006 13960
rect 17313 13957 17325 13960
rect 17359 13988 17371 13991
rect 17402 13988 17408 14000
rect 17359 13960 17408 13988
rect 17359 13957 17371 13960
rect 17313 13951 17371 13957
rect 17402 13948 17408 13960
rect 17460 13988 17466 14000
rect 17880 13988 17908 14028
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 17460 13960 17908 13988
rect 17957 13991 18015 13997
rect 17460 13948 17466 13960
rect 17957 13957 17969 13991
rect 18003 13957 18015 13991
rect 17957 13951 18015 13957
rect 15930 13920 15936 13932
rect 15488 13892 15936 13920
rect 14461 13883 14519 13889
rect 15930 13880 15936 13892
rect 15988 13920 15994 13932
rect 17972 13920 18000 13951
rect 15988 13892 16344 13920
rect 15988 13880 15994 13892
rect 16316 13864 16344 13892
rect 17880 13892 18000 13920
rect 6454 13812 6460 13864
rect 6512 13852 6518 13864
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6512 13824 6561 13852
rect 6512 13812 6518 13824
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8110 13852 8116 13864
rect 7892 13824 8116 13852
rect 7892 13812 7898 13824
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 8478 13852 8484 13864
rect 8439 13824 8484 13852
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 11790 13852 11796 13864
rect 9646 13824 11796 13852
rect 5859 13756 6316 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 9646 13784 9674 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14366 13852 14372 13864
rect 14047 13824 14372 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 9548 13756 9674 13784
rect 9548 13744 9554 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10410 13784 10416 13796
rect 9824 13756 10416 13784
rect 9824 13744 9830 13756
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 12176 13784 12204 13815
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 15304 13824 16160 13852
rect 15304 13784 15332 13824
rect 12176 13756 15332 13784
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 15528 13756 15573 13784
rect 15528 13744 15534 13756
rect 7929 13719 7987 13725
rect 7929 13716 7941 13719
rect 5736 13688 7941 13716
rect 7929 13685 7941 13688
rect 7975 13716 7987 13719
rect 8202 13716 8208 13728
rect 7975 13688 8208 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 10134 13716 10140 13728
rect 8536 13688 10140 13716
rect 8536 13676 8542 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 12618 13716 12624 13728
rect 10551 13688 12624 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 16132 13725 16160 13824
rect 16298 13812 16304 13864
rect 16356 13812 16362 13864
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17402 13852 17408 13864
rect 16960 13824 17408 13852
rect 16758 13784 16764 13796
rect 16592 13756 16764 13784
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 14608 13688 15301 13716
rect 14608 13676 14614 13688
rect 15289 13685 15301 13688
rect 15335 13685 15347 13719
rect 15289 13679 15347 13685
rect 16117 13719 16175 13725
rect 16117 13685 16129 13719
rect 16163 13716 16175 13719
rect 16592 13716 16620 13756
rect 16758 13744 16764 13756
rect 16816 13784 16822 13796
rect 16960 13793 16988 13824
rect 17402 13812 17408 13824
rect 17460 13852 17466 13864
rect 17880 13852 17908 13892
rect 17460 13824 17908 13852
rect 17460 13812 17466 13824
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 16816 13756 16957 13784
rect 16816 13744 16822 13756
rect 16945 13753 16957 13756
rect 16991 13753 17003 13787
rect 16945 13747 17003 13753
rect 18325 13787 18383 13793
rect 18325 13753 18337 13787
rect 18371 13784 18383 13787
rect 18506 13784 18512 13796
rect 18371 13756 18512 13784
rect 18371 13753 18383 13756
rect 18325 13747 18383 13753
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 16163 13688 16620 13716
rect 16163 13685 16175 13688
rect 16117 13679 16175 13685
rect 16666 13676 16672 13728
rect 16724 13716 16730 13728
rect 17957 13719 18015 13725
rect 17957 13716 17969 13719
rect 16724 13688 17969 13716
rect 16724 13676 16730 13688
rect 17957 13685 17969 13688
rect 18003 13685 18015 13719
rect 17957 13679 18015 13685
rect 18230 13676 18236 13728
rect 18288 13716 18294 13728
rect 18690 13716 18696 13728
rect 18288 13688 18696 13716
rect 18288 13676 18294 13688
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 4154 13512 4160 13524
rect 1995 13484 3832 13512
rect 4115 13484 4160 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2133 13447 2191 13453
rect 2133 13413 2145 13447
rect 2179 13444 2191 13447
rect 2590 13444 2596 13456
rect 2179 13416 2596 13444
rect 2179 13413 2191 13416
rect 2133 13407 2191 13413
rect 2590 13404 2596 13416
rect 2648 13404 2654 13456
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13413 2743 13447
rect 3804 13444 3832 13484
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4387 13484 5764 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4801 13447 4859 13453
rect 4801 13444 4813 13447
rect 3804 13416 4813 13444
rect 2685 13407 2743 13413
rect 4801 13413 4813 13416
rect 4847 13413 4859 13447
rect 5736 13444 5764 13484
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5868 13484 5913 13512
rect 5868 13472 5874 13484
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6638 13512 6644 13524
rect 6052 13484 6097 13512
rect 6599 13484 6644 13512
rect 6052 13472 6058 13484
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 6880 13484 7420 13512
rect 6880 13472 6886 13484
rect 5736 13416 7052 13444
rect 4801 13407 4859 13413
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2700 13376 2728 13407
rect 2004 13348 2728 13376
rect 3053 13379 3111 13385
rect 2004 13336 2010 13348
rect 3053 13345 3065 13379
rect 3099 13376 3111 13379
rect 3510 13376 3516 13388
rect 3099 13348 3516 13376
rect 3099 13345 3111 13348
rect 3053 13339 3111 13345
rect 3510 13336 3516 13348
rect 3568 13376 3574 13388
rect 3568 13348 3643 13376
rect 3568 13336 3574 13348
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 3615 13308 3643 13348
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 5684 13348 6500 13376
rect 5684 13336 5690 13348
rect 1627 13280 3556 13308
rect 3615 13280 4109 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 1210 13200 1216 13252
rect 1268 13240 1274 13252
rect 1268 13212 2636 13240
rect 1268 13200 1274 13212
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2608 13181 2636 13212
rect 2593 13175 2651 13181
rect 2593 13141 2605 13175
rect 2639 13141 2651 13175
rect 3528 13172 3556 13280
rect 3970 13240 3976 13252
rect 3931 13212 3976 13240
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4081 13240 4109 13280
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5224 13280 5269 13308
rect 5224 13268 5230 13280
rect 4081 13212 4752 13240
rect 4183 13175 4241 13181
rect 4183 13172 4195 13175
rect 3528 13144 4195 13172
rect 2593 13135 2651 13141
rect 4183 13141 4195 13144
rect 4229 13172 4241 13175
rect 4614 13172 4620 13184
rect 4229 13144 4620 13172
rect 4229 13141 4241 13144
rect 4183 13135 4241 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4724 13172 4752 13212
rect 4890 13200 4896 13252
rect 4948 13240 4954 13252
rect 4985 13243 5043 13249
rect 4985 13240 4997 13243
rect 4948 13212 4997 13240
rect 4948 13200 4954 13212
rect 4985 13209 4997 13212
rect 5031 13209 5043 13243
rect 5629 13243 5687 13249
rect 5629 13240 5641 13243
rect 4985 13203 5043 13209
rect 5276 13212 5641 13240
rect 5276 13172 5304 13212
rect 5629 13209 5641 13212
rect 5675 13240 5687 13243
rect 6178 13240 6184 13252
rect 5675 13212 6184 13240
rect 5675 13209 5687 13212
rect 5629 13203 5687 13209
rect 6178 13200 6184 13212
rect 6236 13200 6242 13252
rect 6472 13249 6500 13348
rect 7024 13308 7052 13416
rect 7392 13376 7420 13484
rect 7466 13472 7472 13524
rect 7524 13472 7530 13524
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 11514 13512 11520 13524
rect 7708 13484 11520 13512
rect 7708 13472 7714 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 11940 13484 14657 13512
rect 11940 13472 11946 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 16942 13512 16948 13524
rect 15335 13484 16948 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17368 13484 17417 13512
rect 17368 13472 17374 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 18325 13515 18383 13521
rect 18325 13481 18337 13515
rect 18371 13512 18383 13515
rect 18690 13512 18696 13524
rect 18371 13484 18696 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 7484 13444 7512 13472
rect 7742 13444 7748 13456
rect 7484 13416 7748 13444
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 8573 13447 8631 13453
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 9490 13444 9496 13456
rect 8619 13416 9496 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 9490 13404 9496 13416
rect 9548 13404 9554 13456
rect 10962 13444 10968 13456
rect 10704 13416 10968 13444
rect 7392 13348 8156 13376
rect 7098 13308 7104 13320
rect 7024 13280 7104 13308
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7742 13308 7748 13320
rect 7703 13280 7748 13308
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13209 6515 13243
rect 6457 13203 6515 13209
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 8128 13240 8156 13348
rect 8202 13336 8208 13388
rect 8260 13376 8266 13388
rect 9398 13376 9404 13388
rect 8260 13348 9404 13376
rect 8260 13336 8266 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 10219 13379 10277 13385
rect 10219 13376 10231 13379
rect 9916 13348 10231 13376
rect 9916 13336 9922 13348
rect 10219 13345 10231 13348
rect 10265 13345 10277 13379
rect 10219 13339 10277 13345
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13376 10563 13379
rect 10704 13376 10732 13416
rect 10962 13404 10968 13416
rect 11020 13404 11026 13456
rect 18138 13444 18144 13456
rect 15580 13416 17264 13444
rect 18099 13416 18144 13444
rect 10551 13348 10732 13376
rect 10781 13379 10839 13385
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 13262 13376 13268 13388
rect 10827 13348 13268 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 13725 13379 13783 13385
rect 13725 13376 13737 13379
rect 13596 13348 13737 13376
rect 13596 13336 13602 13348
rect 13725 13345 13737 13348
rect 13771 13345 13783 13379
rect 13725 13339 13783 13345
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15580 13376 15608 13416
rect 16485 13379 16543 13385
rect 16485 13376 16497 13379
rect 14792 13348 15608 13376
rect 15672 13348 16497 13376
rect 14792 13336 14798 13348
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8570 13308 8576 13320
rect 8435 13280 8576 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8570 13268 8576 13280
rect 8628 13308 8634 13320
rect 9306 13308 9312 13320
rect 8628 13280 9312 13308
rect 8628 13268 8634 13280
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10410 13317 10416 13320
rect 10367 13311 10416 13317
rect 10367 13277 10379 13311
rect 10413 13277 10416 13311
rect 10367 13271 10416 13277
rect 10410 13268 10416 13271
rect 10468 13268 10474 13320
rect 11238 13308 11244 13320
rect 11199 13280 11244 13308
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 8205 13243 8263 13249
rect 8205 13240 8217 13243
rect 7432 13212 7604 13240
rect 8128 13212 8217 13240
rect 7432 13200 7438 13212
rect 4724 13144 5304 13172
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 5829 13175 5887 13181
rect 5829 13172 5841 13175
rect 5408 13144 5841 13172
rect 5408 13132 5414 13144
rect 5829 13141 5841 13144
rect 5875 13141 5887 13175
rect 5829 13135 5887 13141
rect 5994 13132 6000 13184
rect 6052 13172 6058 13184
rect 6657 13175 6715 13181
rect 6657 13172 6669 13175
rect 6052 13144 6669 13172
rect 6052 13132 6058 13144
rect 6657 13141 6669 13144
rect 6703 13141 6715 13175
rect 6657 13135 6715 13141
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13172 6883 13175
rect 7466 13172 7472 13184
rect 6871 13144 7472 13172
rect 6871 13141 6883 13144
rect 6825 13135 6883 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7576 13181 7604 13212
rect 8205 13209 8217 13212
rect 8251 13240 8263 13243
rect 8478 13240 8484 13252
rect 8251 13212 8484 13240
rect 8251 13209 8263 13212
rect 8205 13203 8263 13209
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 7561 13175 7619 13181
rect 7561 13141 7573 13175
rect 7607 13141 7619 13175
rect 9582 13172 9588 13184
rect 9543 13144 9588 13172
rect 7561 13135 7619 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 11440 13172 11468 13271
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11572 13280 11897 13308
rect 11572 13268 11578 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 12894 13308 12900 13320
rect 12855 13280 12900 13308
rect 11885 13271 11943 13277
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15102 13308 15108 13320
rect 14875 13280 15108 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15672 13317 15700 13348
rect 16485 13345 16497 13348
rect 16531 13376 16543 13379
rect 17126 13376 17132 13388
rect 16531 13348 17132 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15344 13280 15485 13308
rect 15344 13268 15350 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15804 13280 16129 13308
rect 15804 13268 15810 13280
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 16117 13271 16175 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16448 13280 16957 13308
rect 16448 13268 16454 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17236 13317 17264 13416
rect 18138 13404 18144 13416
rect 18196 13404 18202 13456
rect 17221 13311 17279 13317
rect 17092 13280 17137 13308
rect 17092 13268 17098 13280
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 15764 13240 15792 13268
rect 15212 13212 15792 13240
rect 15212 13184 15240 13212
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 17184 13212 17877 13240
rect 17184 13200 17190 13212
rect 17865 13209 17877 13212
rect 17911 13209 17923 13243
rect 17865 13203 17923 13209
rect 10008 13144 11468 13172
rect 13081 13175 13139 13181
rect 10008 13132 10014 13144
rect 13081 13141 13093 13175
rect 13127 13172 13139 13175
rect 13354 13172 13360 13184
rect 13127 13144 13360 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 16206 13132 16212 13184
rect 16264 13172 16270 13184
rect 18506 13172 18512 13184
rect 16264 13144 18512 13172
rect 16264 13132 16270 13144
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 1302 12928 1308 12980
rect 1360 12968 1366 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 1360 12940 2145 12968
rect 1360 12928 1366 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 4798 12968 4804 12980
rect 4755 12940 4804 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 7558 12968 7564 12980
rect 5132 12940 7564 12968
rect 5132 12928 5138 12940
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7760 12940 7941 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2682 12900 2688 12912
rect 1995 12872 2688 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 4359 12903 4417 12909
rect 4359 12900 4371 12903
rect 4304 12872 4371 12900
rect 4304 12860 4310 12872
rect 4359 12869 4371 12872
rect 4405 12869 4417 12903
rect 4359 12863 4417 12869
rect 4522 12860 4528 12912
rect 4580 12900 4586 12912
rect 4580 12872 4625 12900
rect 4580 12860 4586 12872
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6794 12903 6852 12909
rect 6794 12900 6806 12903
rect 6512 12872 6806 12900
rect 6512 12860 6518 12872
rect 6794 12869 6806 12872
rect 6840 12869 6852 12903
rect 6794 12863 6852 12869
rect 7760 12900 7788 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 8849 12971 8907 12977
rect 8849 12968 8861 12971
rect 8812 12940 8861 12968
rect 8812 12928 8818 12940
rect 8849 12937 8861 12940
rect 8895 12937 8907 12971
rect 8849 12931 8907 12937
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10284 12940 10333 12968
rect 10284 12928 10290 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 10321 12931 10379 12937
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10928 12940 10977 12968
rect 10928 12928 10934 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11664 12940 11805 12968
rect 11664 12928 11670 12940
rect 11793 12937 11805 12940
rect 11839 12937 11851 12971
rect 11793 12931 11851 12937
rect 12989 12971 13047 12977
rect 12989 12937 13001 12971
rect 13035 12968 13047 12971
rect 13446 12968 13452 12980
rect 13035 12940 13452 12968
rect 13035 12937 13047 12940
rect 12989 12931 13047 12937
rect 7760 12872 11008 12900
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 3697 12835 3755 12841
rect 1627 12804 3648 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3050 12764 3056 12776
rect 3011 12736 3056 12764
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 3510 12764 3516 12776
rect 3471 12736 3516 12764
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3620 12764 3648 12804
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3786 12832 3792 12844
rect 3743 12804 3792 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5920 12832 6132 12836
rect 7760 12832 7788 12872
rect 10980 12844 11008 12872
rect 5675 12808 7788 12832
rect 5675 12804 5948 12808
rect 6104 12804 7788 12808
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8904 12804 9045 12832
rect 8904 12792 8910 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9490 12832 9496 12844
rect 9180 12804 9225 12832
rect 9324 12804 9496 12832
rect 9180 12792 9186 12804
rect 4798 12764 4804 12776
rect 3620 12736 4804 12764
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 3694 12696 3700 12708
rect 3007 12668 3700 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 3804 12668 4568 12696
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 3804 12628 3832 12668
rect 1995 12600 3832 12628
rect 3881 12631 3939 12637
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4338 12628 4344 12640
rect 3927 12600 4344 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4540 12628 4568 12668
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5552 12696 5580 12727
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6144 12736 6561 12764
rect 6144 12724 6150 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 9324 12764 9352 12804
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9640 12804 9873 12832
rect 9640 12792 9646 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10778 12832 10784 12844
rect 10551 12804 10784 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11808 12832 11836 12931
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 17195 12971 17253 12977
rect 17195 12968 17207 12971
rect 13771 12940 17207 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 17195 12937 17207 12940
rect 17241 12937 17253 12971
rect 17862 12968 17868 12980
rect 17823 12940 17868 12968
rect 17195 12931 17253 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18196 12940 18245 12968
rect 18196 12928 18202 12940
rect 18233 12937 18245 12940
rect 18279 12937 18291 12971
rect 18233 12931 18291 12937
rect 18322 12928 18328 12980
rect 18380 12928 18386 12980
rect 13906 12900 13912 12912
rect 13556 12872 13912 12900
rect 13556 12841 13584 12872
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 17402 12900 17408 12912
rect 14792 12872 15700 12900
rect 17363 12872 17408 12900
rect 14792 12860 14798 12872
rect 15672 12844 15700 12872
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 18340 12900 18368 12928
rect 18064 12872 18368 12900
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11808 12804 12265 12832
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 7708 12736 9352 12764
rect 7708 12724 7714 12736
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 11238 12764 11244 12776
rect 9456 12736 11244 12764
rect 9456 12724 9462 12736
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 13096 12764 13124 12795
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14642 12832 14648 12844
rect 14231 12804 14648 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14976 12804 15025 12832
rect 14976 12792 14982 12804
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15013 12795 15071 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 17770 12832 17776 12844
rect 16448 12804 17776 12832
rect 16448 12792 16454 12804
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18064 12841 18092 12872
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 15194 12764 15200 12776
rect 13096 12736 15200 12764
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 18340 12764 18368 12795
rect 16264 12736 18368 12764
rect 16264 12724 16270 12736
rect 5626 12696 5632 12708
rect 4764 12668 5632 12696
rect 4764 12656 4770 12668
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 5997 12699 6055 12705
rect 5997 12665 6009 12699
rect 6043 12696 6055 12699
rect 6454 12696 6460 12708
rect 6043 12668 6460 12696
rect 6043 12665 6055 12668
rect 5997 12659 6055 12665
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 7558 12656 7564 12708
rect 7616 12696 7622 12708
rect 11790 12696 11796 12708
rect 7616 12668 11796 12696
rect 7616 12656 7622 12668
rect 11790 12656 11796 12668
rect 11848 12656 11854 12708
rect 12437 12699 12495 12705
rect 12437 12665 12449 12699
rect 12483 12696 12495 12699
rect 15470 12696 15476 12708
rect 12483 12668 14872 12696
rect 15431 12668 15476 12696
rect 12483 12665 12495 12668
rect 12437 12659 12495 12665
rect 14844 12640 14872 12668
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 16298 12696 16304 12708
rect 16259 12668 16304 12696
rect 16298 12656 16304 12668
rect 16356 12656 16362 12708
rect 17954 12696 17960 12708
rect 17236 12668 17960 12696
rect 6914 12628 6920 12640
rect 4540 12600 6920 12628
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 9398 12628 9404 12640
rect 7524 12600 9404 12628
rect 7524 12588 7530 12600
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 10134 12628 10140 12640
rect 9723 12600 10140 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14056 12600 14381 12628
rect 14056 12588 14062 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 14826 12588 14832 12640
rect 14884 12588 14890 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17236 12637 17264 12668
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 18322 12656 18328 12708
rect 18380 12696 18386 12708
rect 18506 12696 18512 12708
rect 18380 12668 18512 12696
rect 18380 12656 18386 12668
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 16908 12600 17049 12628
rect 16908 12588 16914 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 17221 12631 17279 12637
rect 17221 12597 17233 12631
rect 17267 12597 17279 12631
rect 17221 12591 17279 12597
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 2924 12396 4568 12424
rect 2924 12384 2930 12396
rect 4540 12356 4568 12396
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4985 12427 5043 12433
rect 4985 12424 4997 12427
rect 4672 12396 4997 12424
rect 4672 12384 4678 12396
rect 4985 12393 4997 12396
rect 5031 12393 5043 12427
rect 6546 12424 6552 12436
rect 6507 12396 6552 12424
rect 4985 12387 5043 12393
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 6880 12396 7205 12424
rect 6880 12384 6886 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9088 12396 9229 12424
rect 9088 12384 9094 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9824 12396 9873 12424
rect 9824 12384 9830 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 9861 12387 9919 12393
rect 10689 12427 10747 12433
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 11054 12424 11060 12436
rect 10735 12396 11060 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11790 12424 11796 12436
rect 11751 12396 11796 12424
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 15010 12424 15016 12436
rect 14783 12396 15016 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 16669 12427 16727 12433
rect 15304 12396 16528 12424
rect 5997 12359 6055 12365
rect 4540 12328 5212 12356
rect 934 12248 940 12300
rect 992 12288 998 12300
rect 1302 12288 1308 12300
rect 992 12260 1308 12288
rect 992 12248 998 12260
rect 1302 12248 1308 12260
rect 1360 12248 1366 12300
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1581 12291 1639 12297
rect 1581 12288 1593 12291
rect 1544 12260 1593 12288
rect 1544 12248 1550 12260
rect 1581 12257 1593 12260
rect 1627 12257 1639 12291
rect 1581 12251 1639 12257
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 3844 12260 4476 12288
rect 3844 12248 3850 12260
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 1780 12192 3985 12220
rect 1302 12112 1308 12164
rect 1360 12152 1366 12164
rect 1780 12152 1808 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 1360 12124 1808 12152
rect 1848 12155 1906 12161
rect 1360 12112 1366 12124
rect 1848 12121 1860 12155
rect 1894 12121 1906 12155
rect 1848 12115 1906 12121
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 1872 12084 1900 12115
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 4062 12152 4068 12164
rect 3752 12124 4068 12152
rect 3752 12112 3758 12124
rect 4062 12112 4068 12124
rect 4120 12152 4126 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 4120 12124 4169 12152
rect 4120 12112 4126 12124
rect 4157 12121 4169 12124
rect 4203 12121 4215 12155
rect 4157 12115 4215 12121
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12121 4399 12155
rect 4448 12152 4476 12260
rect 5184 12220 5212 12328
rect 5997 12325 6009 12359
rect 6043 12356 6055 12359
rect 6638 12356 6644 12368
rect 6043 12328 6644 12356
rect 6043 12325 6055 12328
rect 5997 12319 6055 12325
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 6788 12328 8616 12356
rect 6788 12316 6794 12328
rect 8478 12288 8484 12300
rect 8404 12260 8484 12288
rect 5629 12223 5687 12229
rect 5184 12192 5488 12220
rect 4982 12161 4988 12164
rect 4969 12155 4988 12161
rect 4969 12152 4981 12155
rect 4448 12124 4981 12152
rect 4341 12115 4399 12121
rect 4969 12121 4981 12124
rect 4969 12115 4988 12121
rect 2958 12084 2964 12096
rect 1820 12056 1900 12084
rect 2919 12056 2964 12084
rect 1820 12044 1826 12056
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 4356 12084 4384 12115
rect 4982 12112 4988 12115
rect 5040 12112 5046 12164
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 5169 12155 5227 12161
rect 5169 12152 5181 12155
rect 5132 12124 5181 12152
rect 5132 12112 5138 12124
rect 5169 12121 5181 12124
rect 5215 12121 5227 12155
rect 5169 12115 5227 12121
rect 4798 12084 4804 12096
rect 3476 12056 4384 12084
rect 4759 12056 4804 12084
rect 3476 12044 3482 12056
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5460 12084 5488 12192
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5994 12220 6000 12232
rect 5675 12192 6000 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12152 5871 12155
rect 6178 12152 6184 12164
rect 5859 12124 6184 12152
rect 5859 12121 5871 12124
rect 5813 12115 5871 12121
rect 6178 12112 6184 12124
rect 6236 12152 6242 12164
rect 6362 12152 6368 12164
rect 6236 12124 6368 12152
rect 6236 12112 6242 12124
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 6656 12152 6684 12183
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 6880 12192 7113 12220
rect 6880 12180 6886 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7742 12220 7748 12232
rect 7703 12192 7748 12220
rect 7101 12183 7159 12189
rect 7742 12180 7748 12192
rect 7800 12220 7806 12232
rect 8294 12220 8300 12232
rect 7800 12192 8300 12220
rect 7800 12180 7806 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8404 12229 8432 12260
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8588 12288 8616 12328
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 10870 12356 10876 12368
rect 9180 12328 10876 12356
rect 9180 12316 9186 12328
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 13725 12359 13783 12365
rect 13725 12325 13737 12359
rect 13771 12356 13783 12359
rect 15304 12356 15332 12396
rect 13771 12328 15332 12356
rect 15381 12359 15439 12365
rect 13771 12325 13783 12328
rect 13725 12319 13783 12325
rect 15381 12325 15393 12359
rect 15427 12356 15439 12359
rect 16390 12356 16396 12368
rect 15427 12328 16396 12356
rect 15427 12325 15439 12328
rect 15381 12319 15439 12325
rect 16390 12316 16396 12328
rect 16448 12316 16454 12368
rect 16500 12356 16528 12396
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 16942 12424 16948 12436
rect 16715 12396 16948 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17494 12424 17500 12436
rect 17267 12396 17500 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 19242 12356 19248 12368
rect 16500 12328 19248 12356
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 10410 12288 10416 12300
rect 8588 12260 10416 12288
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 12802 12288 12808 12300
rect 10520 12260 12808 12288
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8389 12183 8447 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8996 12192 9413 12220
rect 8996 12180 9002 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 9401 12183 9459 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10520 12229 10548 12260
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 15838 12288 15844 12300
rect 14568 12260 15844 12288
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12189 10563 12223
rect 11146 12220 11152 12232
rect 11107 12192 11152 12220
rect 10505 12183 10563 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 14568 12229 14596 12260
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 16022 12288 16028 12300
rect 15983 12260 16028 12288
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17460 12260 18276 12288
rect 17460 12248 17466 12260
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11296 12192 11989 12220
rect 11296 12180 11302 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 7466 12152 7472 12164
rect 6656 12124 7472 12152
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 12986 12152 12992 12164
rect 7944 12124 12992 12152
rect 7650 12084 7656 12096
rect 5460 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7944 12093 7972 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 13096 12152 13124 12183
rect 15010 12152 15016 12164
rect 13096 12124 15016 12152
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15212 12152 15240 12183
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 16298 12220 16304 12232
rect 15344 12192 16304 12220
rect 15344 12180 15350 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17034 12152 17040 12164
rect 15212 12124 17040 12152
rect 17034 12112 17040 12124
rect 17092 12112 17098 12164
rect 17310 12152 17316 12164
rect 17271 12124 17316 12152
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 17402 12112 17408 12164
rect 17460 12152 17466 12164
rect 18248 12161 18276 12260
rect 18017 12155 18075 12161
rect 18017 12152 18029 12155
rect 17460 12124 18029 12152
rect 17460 12112 17466 12124
rect 18017 12121 18029 12124
rect 18063 12121 18075 12155
rect 18017 12115 18075 12121
rect 18233 12155 18291 12161
rect 18233 12121 18245 12155
rect 18279 12121 18291 12155
rect 18233 12115 18291 12121
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 10686 12084 10692 12096
rect 8619 12056 10692 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 16448 12056 17877 12084
rect 16448 12044 16454 12056
rect 17865 12053 17877 12056
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 4430 11880 4436 11892
rect 2924 11852 4436 11880
rect 2924 11840 2930 11852
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 6546 11880 6552 11892
rect 4580 11852 6552 11880
rect 4580 11840 4586 11852
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7742 11880 7748 11892
rect 6687 11852 7748 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9125 11883 9183 11889
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 9398 11880 9404 11892
rect 9171 11852 9404 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9674 11880 9680 11892
rect 9631 11852 9680 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 10284 11852 10333 11880
rect 10284 11840 10290 11852
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 10321 11843 10379 11849
rect 10410 11840 10416 11892
rect 10468 11880 10474 11892
rect 10870 11880 10876 11892
rect 10468 11852 10732 11880
rect 10831 11852 10876 11880
rect 10468 11840 10474 11852
rect 3510 11812 3516 11824
rect 3423 11784 3516 11812
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1544 11716 1593 11744
rect 1544 11704 1550 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1848 11747 1906 11753
rect 1848 11713 1860 11747
rect 1894 11744 1906 11747
rect 2130 11744 2136 11756
rect 1894 11716 2136 11744
rect 1894 11713 1906 11716
rect 1848 11707 1906 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3436 11753 3464 11784
rect 3510 11772 3516 11784
rect 3568 11812 3574 11824
rect 4982 11812 4988 11824
rect 3568 11784 4988 11812
rect 3568 11772 3574 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 5521 11815 5579 11821
rect 5521 11781 5533 11815
rect 5567 11812 5579 11815
rect 5567 11784 5672 11812
rect 5567 11781 5579 11784
rect 5521 11775 5579 11781
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4706 11744 4712 11756
rect 3835 11716 4712 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11676 3571 11679
rect 3602 11676 3608 11688
rect 3559 11648 3608 11676
rect 3559 11645 3571 11648
rect 3513 11639 3571 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 3712 11676 3740 11707
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5258 11744 5264 11756
rect 4948 11716 5264 11744
rect 4948 11704 4954 11716
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5644 11744 5672 11784
rect 5718 11772 5724 11824
rect 5776 11812 5782 11824
rect 5776 11784 5821 11812
rect 5776 11772 5782 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 9490 11812 9496 11824
rect 7708 11784 9496 11812
rect 7708 11772 7714 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 10594 11812 10600 11824
rect 9784 11784 10600 11812
rect 6454 11744 6460 11756
rect 5644 11716 6460 11744
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 7064 11716 7113 11744
rect 7064 11704 7070 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 7926 11744 7932 11756
rect 7883 11716 7932 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9784 11753 9812 11784
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 10704 11812 10732 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14148 11852 14289 11880
rect 14148 11840 14154 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11880 14979 11883
rect 15470 11880 15476 11892
rect 14967 11852 15476 11880
rect 14967 11849 14979 11852
rect 14921 11843 14979 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 17402 11880 17408 11892
rect 15703 11852 17408 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17954 11880 17960 11892
rect 17915 11852 17960 11880
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 19426 11880 19432 11892
rect 18064 11852 19432 11880
rect 10704 11784 11100 11812
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8720 11716 8953 11744
rect 8720 11704 8726 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10870 11744 10876 11756
rect 10831 11716 10876 11744
rect 10229 11707 10287 11713
rect 3878 11676 3884 11688
rect 3712 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4019 11648 4752 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 842 11568 848 11620
rect 900 11608 906 11620
rect 1118 11608 1124 11620
rect 900 11580 1124 11608
rect 900 11568 906 11580
rect 1118 11568 1124 11580
rect 1176 11568 1182 11620
rect 4172 11580 4568 11608
rect 2961 11543 3019 11549
rect 2961 11509 2973 11543
rect 3007 11540 3019 11543
rect 3418 11540 3424 11552
rect 3007 11512 3424 11540
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 3418 11500 3424 11512
rect 3476 11540 3482 11552
rect 4062 11540 4068 11552
rect 3476 11512 4068 11540
rect 3476 11500 3482 11512
rect 4062 11500 4068 11512
rect 4120 11540 4126 11552
rect 4172 11540 4200 11580
rect 4120 11512 4200 11540
rect 4120 11500 4126 11512
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4304 11512 4445 11540
rect 4304 11500 4310 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 4540 11540 4568 11580
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4540 11512 4629 11540
rect 4433 11503 4491 11509
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4724 11540 4752 11648
rect 5074 11636 5080 11688
rect 5132 11676 5138 11688
rect 7282 11676 7288 11688
rect 5132 11648 7288 11676
rect 5132 11636 5138 11648
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 10244 11676 10272 11707
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11072 11753 11100 11784
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 18064 11812 18092 11852
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 18322 11812 18328 11824
rect 15068 11784 18092 11812
rect 18283 11784 18328 11812
rect 15068 11772 15074 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11713 11115 11747
rect 11698 11744 11704 11756
rect 11659 11716 11704 11744
rect 11057 11707 11115 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 13722 11744 13728 11756
rect 13683 11716 13728 11744
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14642 11744 14648 11756
rect 14415 11716 14648 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14826 11744 14832 11756
rect 14787 11716 14832 11744
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 15344 11716 15485 11744
rect 15344 11704 15350 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 9140 11648 10272 11676
rect 13081 11679 13139 11685
rect 5350 11608 5356 11620
rect 5311 11580 5356 11608
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 9140 11608 9168 11648
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 14734 11676 14740 11688
rect 13127 11648 14740 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15672 11676 15700 11707
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 15988 11716 16313 11744
rect 15988 11704 15994 11716
rect 16301 11713 16313 11716
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 18012 11716 18153 11744
rect 18012 11704 18018 11716
rect 18141 11713 18153 11716
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18046 11676 18052 11688
rect 15672 11648 18052 11676
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 7984 11580 9168 11608
rect 7984 11568 7990 11580
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 11422 11608 11428 11620
rect 9456 11580 11428 11608
rect 9456 11568 9462 11580
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 17494 11608 17500 11620
rect 17455 11580 17500 11608
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 5074 11540 5080 11552
rect 4724 11512 5080 11540
rect 4617 11503 4675 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5537 11543 5595 11549
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 5718 11540 5724 11552
rect 5583 11512 5724 11540
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 10870 11540 10876 11552
rect 6328 11512 10876 11540
rect 6328 11500 6334 11512
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 1118 11296 1124 11348
rect 1176 11336 1182 11348
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 1176 11308 3985 11336
rect 1176 11296 1182 11308
rect 3973 11305 3985 11308
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 5258 11336 5264 11348
rect 4203 11308 5264 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 7524 11308 9137 11336
rect 7524 11296 7530 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 9769 11339 9827 11345
rect 9769 11336 9781 11339
rect 9732 11308 9781 11336
rect 9732 11296 9738 11308
rect 9769 11305 9781 11308
rect 9815 11305 9827 11339
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 9769 11299 9827 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 15105 11339 15163 11345
rect 15105 11336 15117 11339
rect 14240 11308 15117 11336
rect 14240 11296 14246 11308
rect 15105 11305 15117 11308
rect 15151 11305 15163 11339
rect 15105 11299 15163 11305
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16172 11308 16221 11336
rect 16172 11296 16178 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 17037 11339 17095 11345
rect 17037 11305 17049 11339
rect 17083 11336 17095 11339
rect 17126 11336 17132 11348
rect 17083 11308 17132 11336
rect 17083 11305 17095 11308
rect 17037 11299 17095 11305
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17368 11308 17509 11336
rect 17368 11296 17374 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 3510 11268 3516 11280
rect 3007 11240 3516 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 5166 11268 5172 11280
rect 4396 11240 5172 11268
rect 4396 11228 4402 11240
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 5350 11228 5356 11280
rect 5408 11268 5414 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 5408 11240 7941 11268
rect 5408 11228 5414 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 7929 11231 7987 11237
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 11054 11268 11060 11280
rect 8168 11240 9444 11268
rect 11015 11240 11060 11268
rect 8168 11228 8174 11240
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1581 11203 1639 11209
rect 1581 11200 1593 11203
rect 1544 11172 1593 11200
rect 1544 11160 1550 11172
rect 1581 11169 1593 11172
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 2924 11172 5856 11200
rect 2924 11160 2930 11172
rect 4522 11132 4528 11144
rect 4483 11104 4528 11132
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5074 11132 5080 11144
rect 5031 11104 5080 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 5224 11104 5273 11132
rect 5224 11092 5230 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5828 11132 5856 11172
rect 5902 11160 5908 11212
rect 5960 11200 5966 11212
rect 6178 11200 6184 11212
rect 5960 11172 6184 11200
rect 5960 11160 5966 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6656 11172 8248 11200
rect 6656 11144 6684 11172
rect 6089 11135 6147 11141
rect 5828 11104 6040 11132
rect 5261 11095 5319 11101
rect 1854 11073 1860 11076
rect 1848 11027 1860 11073
rect 1912 11064 1918 11076
rect 1912 11036 1948 11064
rect 1854 11024 1860 11027
rect 1912 11024 1918 11036
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 2556 11036 5457 11064
rect 2556 11024 2562 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5902 11064 5908 11076
rect 5863 11036 5908 11064
rect 5445 11027 5503 11033
rect 5902 11024 5908 11036
rect 5960 11024 5966 11076
rect 6012 11064 6040 11104
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6270 11132 6276 11144
rect 6135 11104 6276 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6638 11132 6644 11144
rect 6599 11104 6644 11132
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 8110 11132 8116 11144
rect 7208 11104 8116 11132
rect 6730 11064 6736 11076
rect 6012 11036 6736 11064
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 2682 10956 2688 11008
rect 2740 10996 2746 11008
rect 4157 10999 4215 11005
rect 4157 10996 4169 10999
rect 2740 10968 4169 10996
rect 2740 10956 2746 10968
rect 4157 10965 4169 10968
rect 4203 10965 4215 10999
rect 5074 10996 5080 11008
rect 5035 10968 5080 10996
rect 4157 10959 4215 10965
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 7208 10996 7236 11104
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8220 11064 8248 11172
rect 9306 11132 9312 11144
rect 9267 11104 9312 11132
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9416 11132 9444 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 14458 11268 14464 11280
rect 14419 11240 14464 11268
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 14976 11240 15669 11268
rect 14976 11228 14982 11240
rect 15657 11237 15669 11240
rect 15703 11237 15715 11271
rect 15657 11231 15715 11237
rect 17678 11228 17684 11280
rect 17736 11228 17742 11280
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 9548 11172 10425 11200
rect 9548 11160 9554 11172
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 17126 11200 17132 11212
rect 10413 11163 10471 11169
rect 16868 11172 17132 11200
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9416 11104 9965 11132
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 16390 11132 16396 11144
rect 16351 11104 16396 11132
rect 15749 11095 15807 11101
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 8220 11036 11713 11064
rect 11701 11033 11713 11036
rect 11747 11033 11759 11067
rect 15764 11064 15792 11095
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16868 11141 16896 11172
rect 17126 11160 17132 11172
rect 17184 11200 17190 11212
rect 17696 11200 17724 11228
rect 17184 11172 17724 11200
rect 17184 11160 17190 11172
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 16853 11095 16911 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 17920 11104 18337 11132
rect 17920 11092 17926 11104
rect 18325 11101 18337 11104
rect 18371 11132 18383 11135
rect 18506 11132 18512 11144
rect 18371 11104 18512 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 17402 11064 17408 11076
rect 15764 11036 17408 11064
rect 11701 11027 11759 11033
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 5224 10968 7236 10996
rect 5224 10956 5230 10968
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 13320 10968 18153 10996
rect 13320 10956 13326 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 6914 10792 6920 10804
rect 2280 10764 5396 10792
rect 6875 10764 6920 10792
rect 2280 10752 2286 10764
rect 2958 10724 2964 10736
rect 2148 10696 2964 10724
rect 2148 10665 2176 10696
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 5368 10724 5396 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 9309 10795 9367 10801
rect 9309 10761 9321 10795
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10318 10792 10324 10804
rect 10091 10764 10324 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 9324 10724 9352 10755
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15102 10792 15108 10804
rect 15059 10764 15108 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17276 10764 17509 10792
rect 17276 10752 17282 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 18414 10724 18420 10736
rect 3344 10696 5304 10724
rect 5368 10696 9352 10724
rect 17696 10696 18420 10724
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2501 10659 2559 10665
rect 2501 10656 2513 10659
rect 2133 10619 2191 10625
rect 2240 10628 2513 10656
rect 2038 10588 2044 10600
rect 1999 10560 2044 10588
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 2240 10520 2268 10628
rect 2501 10625 2513 10628
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2682 10616 2688 10668
rect 2740 10656 2746 10668
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2740 10628 2881 10656
rect 2740 10616 2746 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 2409 10591 2467 10597
rect 2409 10588 2421 10591
rect 1636 10492 2268 10520
rect 2332 10560 2421 10588
rect 1636 10480 1642 10492
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2332 10452 2360 10560
rect 2409 10557 2421 10560
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 3344 10520 3372 10696
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 3436 10588 3464 10619
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3970 10656 3976 10668
rect 3844 10628 3976 10656
rect 3844 10616 3850 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5276 10665 5304 10696
rect 5005 10659 5063 10665
rect 5005 10656 5017 10659
rect 4580 10628 5017 10656
rect 4580 10616 4586 10628
rect 5005 10625 5017 10628
rect 5051 10625 5063 10659
rect 5005 10619 5063 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 3436 10560 3924 10588
rect 3896 10529 3924 10560
rect 2424 10492 3372 10520
rect 3881 10523 3939 10529
rect 2424 10464 2452 10492
rect 3881 10489 3893 10523
rect 3927 10489 3939 10523
rect 5276 10520 5304 10619
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5905 10659 5963 10665
rect 5905 10656 5917 10659
rect 5592 10628 5917 10656
rect 5592 10616 5598 10628
rect 5905 10625 5917 10628
rect 5951 10625 5963 10659
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 5905 10619 5963 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 7374 10656 7380 10668
rect 7335 10628 7380 10656
rect 6733 10619 6791 10625
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 6748 10588 6776 10619
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9272 10628 9505 10656
rect 9272 10616 9278 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9640 10628 9965 10656
rect 9640 10616 9646 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 15746 10656 15752 10668
rect 15703 10628 15752 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16850 10656 16856 10668
rect 16811 10628 16856 10656
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17696 10665 17724 10696
rect 18414 10684 18420 10696
rect 18472 10684 18478 10736
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 18322 10656 18328 10668
rect 18283 10628 18328 10656
rect 17681 10619 17739 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 5408 10560 6776 10588
rect 5408 10548 5414 10560
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7340 10560 8033 10588
rect 7340 10548 7346 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 8168 10560 10609 10588
rect 8168 10548 8174 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 18598 10588 18604 10600
rect 16347 10560 18604 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 5902 10520 5908 10532
rect 5276 10492 5908 10520
rect 3881 10483 3939 10489
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 17037 10523 17095 10529
rect 17037 10489 17049 10523
rect 17083 10520 17095 10523
rect 18230 10520 18236 10532
rect 17083 10492 18236 10520
rect 17083 10489 17095 10492
rect 17037 10483 17095 10489
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 2280 10424 2360 10452
rect 2280 10412 2286 10424
rect 2406 10412 2412 10464
rect 2464 10412 2470 10464
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 2648 10424 5733 10452
rect 2648 10412 2654 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 4522 10248 4528 10260
rect 2832 10220 4528 10248
rect 2832 10208 2838 10220
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5074 10248 5080 10260
rect 4663 10220 5080 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5258 10208 5264 10260
rect 5316 10248 5322 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5316 10220 5457 10248
rect 5316 10208 5322 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6546 10248 6552 10260
rect 5592 10220 6552 10248
rect 5592 10208 5598 10220
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 8076 10220 8125 10248
rect 8076 10208 8082 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 8113 10211 8171 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9769 10251 9827 10257
rect 9769 10248 9781 10251
rect 9364 10220 9781 10248
rect 9364 10208 9370 10220
rect 9769 10217 9781 10220
rect 9815 10217 9827 10251
rect 9769 10211 9827 10217
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 15436 10220 15669 10248
rect 15436 10208 15442 10220
rect 2746 10152 9352 10180
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1544 10084 1593 10112
rect 1544 10072 1550 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1596 10044 1624 10075
rect 2406 10044 2412 10056
rect 1596 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 1848 9979 1906 9985
rect 1848 9945 1860 9979
rect 1894 9976 1906 9979
rect 2222 9976 2228 9988
rect 1894 9948 2228 9976
rect 1894 9945 1906 9948
rect 1848 9939 1906 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 2746 9908 2774 10152
rect 2958 10072 2964 10124
rect 3016 10072 3022 10124
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3108 10084 4109 10112
rect 3108 10072 3114 10084
rect 2976 9976 3004 10072
rect 4081 10053 4109 10084
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 7469 10115 7527 10121
rect 7469 10112 7481 10115
rect 5132 10084 7481 10112
rect 5132 10072 5138 10084
rect 7469 10081 7481 10084
rect 7515 10081 7527 10115
rect 7469 10075 7527 10081
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4066 10047 4124 10053
rect 4066 10013 4078 10047
rect 4112 10013 4124 10047
rect 4246 10044 4252 10056
rect 4207 10016 4252 10044
rect 4066 10007 4124 10013
rect 3050 9976 3056 9988
rect 2976 9948 3056 9976
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 2004 9880 2774 9908
rect 2961 9911 3019 9917
rect 2004 9868 2010 9880
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3418 9908 3424 9920
rect 3007 9880 3424 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3418 9868 3424 9880
rect 3476 9908 3482 9920
rect 3786 9908 3792 9920
rect 3476 9880 3792 9908
rect 3476 9868 3482 9880
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 3988 9908 4016 10007
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4479 10047 4537 10053
rect 4479 10013 4491 10047
rect 4525 10044 4537 10047
rect 4706 10044 4712 10056
rect 4525 10016 4712 10044
rect 4525 10013 4537 10016
rect 4479 10007 4537 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 5040 10016 5273 10044
rect 5040 10004 5046 10016
rect 5261 10013 5273 10016
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 4154 9936 4160 9988
rect 4212 9976 4218 9988
rect 4341 9979 4399 9985
rect 4341 9976 4353 9979
rect 4212 9948 4353 9976
rect 4212 9936 4218 9948
rect 4341 9945 4353 9948
rect 4387 9945 4399 9979
rect 4341 9939 4399 9945
rect 5077 9979 5135 9985
rect 5077 9945 5089 9979
rect 5123 9976 5135 9979
rect 5442 9976 5448 9988
rect 5123 9948 5448 9976
rect 5123 9945 5135 9948
rect 5077 9939 5135 9945
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 6288 9976 6316 10007
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6696 10016 7389 10044
rect 6696 10004 6702 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7377 10007 7435 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8018 10044 8024 10056
rect 7979 10016 8024 10044
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 9324 10053 9352 10152
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9674 10044 9680 10056
rect 9355 10016 9680 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 15488 10044 15516 10220
rect 15657 10217 15669 10220
rect 15703 10217 15715 10251
rect 15657 10211 15715 10217
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 16264 10220 16313 10248
rect 16264 10208 16270 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 17402 10248 17408 10260
rect 17363 10220 17408 10248
rect 16301 10211 16359 10217
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 16761 10183 16819 10189
rect 16761 10180 16773 10183
rect 15620 10152 16773 10180
rect 15620 10140 15626 10152
rect 16761 10149 16773 10152
rect 16807 10149 16819 10183
rect 16761 10143 16819 10149
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 15488 10016 16957 10044
rect 16945 10013 16957 10016
rect 16991 10013 17003 10047
rect 17586 10044 17592 10056
rect 17547 10016 17592 10044
rect 16945 10007 17003 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 10502 9976 10508 9988
rect 6288 9948 10508 9976
rect 10502 9936 10508 9948
rect 10560 9936 10566 9988
rect 4430 9908 4436 9920
rect 3988 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5258 9908 5264 9920
rect 4672 9880 5264 9908
rect 4672 9868 4678 9880
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6086 9908 6092 9920
rect 6047 9880 6092 9908
rect 6086 9868 6092 9880
rect 6144 9868 6150 9920
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2924 9676 5856 9704
rect 2924 9664 2930 9676
rect 2406 9636 2412 9648
rect 1596 9608 2412 9636
rect 1596 9577 1624 9608
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 3697 9639 3755 9645
rect 3697 9636 3709 9639
rect 2648 9608 3709 9636
rect 2648 9596 2654 9608
rect 3697 9605 3709 9608
rect 3743 9636 3755 9639
rect 3743 9608 3924 9636
rect 3743 9605 3755 9608
rect 3697 9599 3755 9605
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 1848 9571 1906 9577
rect 1848 9537 1860 9571
rect 1894 9568 1906 9571
rect 3421 9571 3479 9577
rect 1894 9540 2728 9568
rect 1894 9537 1906 9540
rect 1848 9531 1906 9537
rect 2700 9364 2728 9540
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3510 9568 3516 9580
rect 3467 9540 3516 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3786 9568 3792 9580
rect 3660 9540 3705 9568
rect 3747 9540 3792 9568
rect 3660 9528 3666 9540
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3896 9500 3924 9608
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4614 9636 4620 9648
rect 4212 9608 4620 9636
rect 4212 9596 4218 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4890 9636 4896 9648
rect 4851 9608 4896 9636
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5718 9636 5724 9648
rect 5679 9608 5724 9636
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 5828 9636 5856 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 7558 9704 7564 9716
rect 5960 9676 7564 9704
rect 5960 9664 5966 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7837 9707 7895 9713
rect 7837 9673 7849 9707
rect 7883 9673 7895 9707
rect 17678 9704 17684 9716
rect 7837 9667 7895 9673
rect 16316 9676 17684 9704
rect 7852 9636 7880 9667
rect 5828 9608 7880 9636
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 16316 9645 16344 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 9769 9639 9827 9645
rect 9769 9636 9781 9639
rect 9732 9608 9781 9636
rect 9732 9596 9738 9608
rect 9769 9605 9781 9608
rect 9815 9605 9827 9639
rect 9769 9599 9827 9605
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9605 16359 9639
rect 17954 9636 17960 9648
rect 16301 9599 16359 9605
rect 17696 9608 17960 9636
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 5350 9568 5356 9580
rect 4120 9540 4844 9568
rect 5311 9540 5356 9568
rect 4120 9528 4126 9540
rect 4154 9500 4160 9512
rect 2832 9472 3004 9500
rect 3896 9472 4160 9500
rect 2832 9460 2838 9472
rect 2976 9441 3004 9472
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4430 9500 4436 9512
rect 4391 9472 4436 9500
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 2961 9435 3019 9441
rect 2961 9401 2973 9435
rect 3007 9432 3019 9435
rect 3878 9432 3884 9444
rect 3007 9404 3884 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 3973 9435 4031 9441
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 4338 9432 4344 9444
rect 4019 9404 4344 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 4614 9432 4620 9444
rect 4575 9404 4620 9432
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 4816 9432 4844 9540
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5500 9540 5549 9568
rect 5500 9528 5506 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8202 9568 8208 9580
rect 8067 9540 8208 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 6748 9500 6776 9531
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9122 9568 9128 9580
rect 9083 9540 9128 9568
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 17696 9577 17724 9608
rect 17954 9596 17960 9608
rect 18012 9636 18018 9648
rect 19058 9636 19064 9648
rect 18012 9608 19064 9636
rect 18012 9596 18018 9608
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9568 15807 9571
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 15795 9540 17049 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 17037 9537 17049 9540
rect 17083 9568 17095 9571
rect 17681 9571 17739 9577
rect 17083 9540 17632 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 5040 9472 6776 9500
rect 5040 9460 5046 9472
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 17604 9500 17632 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 18322 9568 18328 9580
rect 18283 9540 18328 9568
rect 17681 9531 17739 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 19150 9500 19156 9512
rect 15252 9472 17540 9500
rect 17604 9472 19156 9500
rect 15252 9460 15258 9472
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 4816 9404 7205 9432
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 14642 9392 14648 9444
rect 14700 9432 14706 9444
rect 17512 9441 17540 9472
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 14700 9404 16865 9432
rect 14700 9392 14706 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16853 9395 16911 9401
rect 17497 9435 17555 9441
rect 17497 9401 17509 9435
rect 17543 9401 17555 9435
rect 17497 9395 17555 9401
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 2700 9336 6561 9364
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 6549 9327 6607 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 4982 9160 4988 9172
rect 2372 9132 4988 9160
rect 2372 9120 2378 9132
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7064 9132 7481 9160
rect 7064 9120 7070 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 8110 9160 8116 9172
rect 8071 9132 8116 9160
rect 7469 9123 7527 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 9125 9163 9183 9169
rect 9125 9160 9137 9163
rect 8720 9132 9137 9160
rect 8720 9120 8726 9132
rect 9125 9129 9137 9132
rect 9171 9129 9183 9163
rect 17126 9160 17132 9172
rect 17087 9132 17132 9160
rect 9125 9123 9183 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 18322 9160 18328 9172
rect 18283 9132 18328 9160
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 3694 9052 3700 9104
rect 3752 9092 3758 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 3752 9064 4077 9092
rect 3752 9052 3758 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 4065 9055 4123 9061
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 4893 9095 4951 9101
rect 4893 9092 4905 9095
rect 4580 9064 4905 9092
rect 4580 9052 4586 9064
rect 4893 9061 4905 9064
rect 4939 9061 4951 9095
rect 4893 9055 4951 9061
rect 6365 9095 6423 9101
rect 6365 9061 6377 9095
rect 6411 9092 6423 9095
rect 8018 9092 8024 9104
rect 6411 9064 8024 9092
rect 6411 9061 6423 9064
rect 6365 9055 6423 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 16669 9095 16727 9101
rect 16669 9061 16681 9095
rect 16715 9092 16727 9095
rect 17862 9092 17868 9104
rect 16715 9064 17868 9092
rect 16715 9061 16727 9064
rect 16669 9055 16727 9061
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 5442 9024 5448 9036
rect 3108 8996 5448 9024
rect 3108 8984 3114 8996
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8925 3019 8959
rect 2961 8919 3019 8925
rect 1946 8888 1952 8900
rect 1596 8860 1952 8888
rect 1596 8829 1624 8860
rect 1946 8848 1952 8860
rect 2004 8888 2010 8900
rect 2590 8888 2596 8900
rect 2004 8860 2596 8888
rect 2004 8848 2010 8860
rect 2590 8848 2596 8860
rect 2648 8848 2654 8900
rect 2716 8891 2774 8897
rect 2716 8857 2728 8891
rect 2762 8888 2774 8891
rect 2866 8888 2872 8900
rect 2762 8860 2872 8888
rect 2762 8857 2774 8860
rect 2716 8851 2774 8857
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2976 8820 3004 8919
rect 3436 8900 3464 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 9024 16175 9027
rect 17954 9024 17960 9036
rect 16163 8996 17960 9024
rect 16163 8993 16175 8996
rect 16117 8987 16175 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4798 8956 4804 8968
rect 4212 8928 4804 8956
rect 4212 8916 4218 8928
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 5350 8956 5356 8968
rect 4856 8928 5356 8956
rect 4856 8916 4862 8928
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 6178 8956 6184 8968
rect 6139 8928 6184 8956
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8956 7067 8959
rect 7098 8956 7104 8968
rect 7055 8928 7104 8956
rect 7055 8925 7067 8928
rect 7009 8919 7067 8925
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 3418 8848 3424 8900
rect 3476 8848 3482 8900
rect 4246 8848 4252 8900
rect 4304 8888 4310 8900
rect 4433 8891 4491 8897
rect 4433 8888 4445 8891
rect 4304 8860 4445 8888
rect 4304 8848 4310 8860
rect 4433 8857 4445 8860
rect 4479 8857 4491 8891
rect 4433 8851 4491 8857
rect 4614 8848 4620 8900
rect 4672 8888 4678 8900
rect 5902 8888 5908 8900
rect 4672 8860 5908 8888
rect 4672 8848 4678 8860
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 2464 8792 3004 8820
rect 2464 8780 2470 8792
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3936 8792 3985 8820
rect 3936 8780 3942 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2314 8616 2320 8628
rect 2179 8588 2320 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2464 8588 2973 8616
rect 2464 8576 2470 8588
rect 2961 8585 2973 8588
rect 3007 8616 3019 8619
rect 3326 8616 3332 8628
rect 3007 8588 3332 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3881 8619 3939 8625
rect 3436 8588 3648 8616
rect 1670 8508 1676 8560
rect 1728 8548 1734 8560
rect 1949 8551 2007 8557
rect 1949 8548 1961 8551
rect 1728 8520 1961 8548
rect 1728 8508 1734 8520
rect 1949 8517 1961 8520
rect 1995 8548 2007 8551
rect 2682 8548 2688 8560
rect 1995 8520 2688 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 2682 8508 2688 8520
rect 2740 8548 2746 8560
rect 3436 8548 3464 8588
rect 2740 8520 3464 8548
rect 3513 8551 3571 8557
rect 2740 8508 2746 8520
rect 3513 8517 3525 8551
rect 3559 8517 3571 8551
rect 3513 8511 3571 8517
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 2590 8480 2596 8492
rect 1627 8452 2596 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2774 8480 2780 8492
rect 2735 8452 2780 8480
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3068 8412 3096 8443
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3528 8480 3556 8511
rect 3476 8452 3556 8480
rect 3476 8440 3482 8452
rect 2740 8384 3096 8412
rect 3620 8412 3648 8588
rect 3881 8585 3893 8619
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 7926 8616 7932 8628
rect 4571 8588 7932 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 3718 8551 3776 8557
rect 3718 8517 3730 8551
rect 3764 8548 3776 8551
rect 3896 8548 3924 8579
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 17586 8616 17592 8628
rect 17359 8588 17592 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 3764 8520 3832 8548
rect 3896 8520 5028 8548
rect 3764 8517 3776 8520
rect 3718 8511 3776 8517
rect 3804 8480 3832 8520
rect 4154 8480 4160 8492
rect 3804 8452 4160 8480
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4338 8480 4344 8492
rect 4299 8452 4344 8480
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5000 8489 5028 8520
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5776 8452 5825 8480
rect 5776 8440 5782 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 7190 8480 7196 8492
rect 7151 8452 7196 8480
rect 6733 8443 6791 8449
rect 3694 8412 3700 8424
rect 3620 8384 3700 8412
rect 2740 8372 2746 8384
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 1964 8316 2605 8344
rect 1964 8285 1992 8316
rect 2593 8313 2605 8316
rect 2639 8313 2651 8347
rect 3068 8344 3096 8384
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 6748 8412 6776 8443
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19150 8480 19156 8492
rect 18371 8452 19156 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 4120 8384 7849 8412
rect 4120 8372 4126 8384
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 7837 8375 7895 8381
rect 3068 8316 4384 8344
rect 2593 8307 2651 8313
rect 1949 8279 2007 8285
rect 1949 8245 1961 8279
rect 1995 8245 2007 8279
rect 1949 8239 2007 8245
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 3418 8276 3424 8288
rect 2372 8248 3424 8276
rect 2372 8236 2378 8248
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 3694 8276 3700 8288
rect 3655 8248 3700 8276
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4356 8276 4384 8316
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 4488 8316 6561 8344
rect 4488 8304 4494 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 4614 8276 4620 8288
rect 4356 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5626 8276 5632 8288
rect 5587 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2590 8072 2596 8084
rect 2551 8044 2596 8072
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2740 8044 2789 8072
rect 2740 8032 2746 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 3970 8072 3976 8084
rect 3931 8044 3976 8072
rect 2777 8035 2835 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4706 8072 4712 8084
rect 4667 8044 4712 8072
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 9582 8072 9588 8084
rect 6779 8044 9588 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 3786 8004 3792 8016
rect 1780 7976 3792 8004
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1780 7877 1808 7976
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 7193 8007 7251 8013
rect 7193 8004 7205 8007
rect 6604 7976 7205 8004
rect 6604 7964 6610 7976
rect 7193 7973 7205 7976
rect 7239 7973 7251 8007
rect 7193 7967 7251 7973
rect 5626 7936 5632 7948
rect 2332 7908 3096 7936
rect 2332 7880 2360 7908
rect 3068 7880 3096 7908
rect 4816 7908 5632 7936
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1636 7840 1777 7868
rect 1636 7828 1642 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 1946 7868 1952 7880
rect 1903 7840 1952 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 2314 7868 2320 7880
rect 2179 7840 2320 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 3050 7828 3056 7880
rect 3108 7828 3114 7880
rect 4816 7877 4844 7908
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 4801 7831 4859 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7098 7868 7104 7880
rect 6595 7840 7104 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 2774 7809 2780 7812
rect 2761 7803 2780 7809
rect 2761 7769 2773 7803
rect 2761 7763 2780 7769
rect 2774 7760 2780 7763
rect 2832 7760 2838 7812
rect 2961 7803 3019 7809
rect 2961 7769 2973 7803
rect 3007 7769 3019 7803
rect 2961 7763 3019 7769
rect 566 7692 572 7744
rect 624 7732 630 7744
rect 2314 7732 2320 7744
rect 624 7704 2320 7732
rect 624 7692 630 7704
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2976 7732 3004 7763
rect 2464 7704 3004 7732
rect 2464 7692 2470 7704
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 2188 7500 2421 7528
rect 2188 7488 2194 7500
rect 2409 7497 2421 7500
rect 2455 7497 2467 7531
rect 2409 7491 2467 7497
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3053 7531 3111 7537
rect 3053 7528 3065 7531
rect 2924 7500 3065 7528
rect 2924 7488 2930 7500
rect 3053 7497 3065 7500
rect 3099 7497 3111 7531
rect 5074 7528 5080 7540
rect 3053 7491 3111 7497
rect 4264 7500 5080 7528
rect 1581 7463 1639 7469
rect 1581 7429 1593 7463
rect 1627 7460 1639 7463
rect 1670 7460 1676 7472
rect 1627 7432 1676 7460
rect 1627 7429 1639 7432
rect 1581 7423 1639 7429
rect 1670 7420 1676 7432
rect 1728 7420 1734 7472
rect 1797 7463 1855 7469
rect 1797 7429 1809 7463
rect 1843 7460 1855 7463
rect 4264 7460 4292 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 5810 7528 5816 7540
rect 5675 7500 5816 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6236 7500 6561 7528
rect 6236 7488 6242 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 6549 7491 6607 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 5994 7460 6000 7472
rect 1843 7432 4292 7460
rect 4356 7432 6000 7460
rect 1843 7429 1855 7432
rect 1797 7423 1855 7429
rect 4356 7401 4384 7432
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 1964 7364 2605 7392
rect 934 7216 940 7268
rect 992 7256 998 7268
rect 1964 7265 1992 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2593 7355 2651 7361
rect 2746 7364 3249 7392
rect 2746 7324 2774 7364
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 5810 7392 5816 7404
rect 4571 7364 5672 7392
rect 5771 7364 5816 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 2056 7296 2774 7324
rect 1949 7259 2007 7265
rect 992 7228 1900 7256
rect 992 7216 998 7228
rect 1302 7148 1308 7200
rect 1360 7188 1366 7200
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 1360 7160 1777 7188
rect 1360 7148 1366 7160
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 1872 7188 1900 7228
rect 1949 7225 1961 7259
rect 1995 7225 2007 7259
rect 1949 7219 2007 7225
rect 2056 7188 2084 7296
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3200 7296 3709 7324
rect 3200 7284 3206 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 3697 7287 3755 7293
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4120 7296 4997 7324
rect 4120 7284 4126 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 5644 7324 5672 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 18322 7392 18328 7404
rect 18283 7364 18328 7392
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 6362 7324 6368 7336
rect 5644 7296 6368 7324
rect 4985 7287 5043 7293
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 5902 7256 5908 7268
rect 2372 7228 5908 7256
rect 2372 7216 2378 7228
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 1872 7160 2084 7188
rect 4433 7191 4491 7197
rect 1765 7151 1823 7157
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 6270 7188 6276 7200
rect 4479 7160 6276 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 5997 6987 6055 6993
rect 5997 6984 6009 6987
rect 5868 6956 6009 6984
rect 5868 6944 5874 6956
rect 5997 6953 6009 6956
rect 6043 6953 6055 6987
rect 5997 6947 6055 6953
rect 4154 6916 4160 6928
rect 3988 6888 4160 6916
rect 3878 6848 3884 6860
rect 2746 6820 3884 6848
rect 1118 6740 1124 6792
rect 1176 6780 1182 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1176 6752 1593 6780
rect 1176 6740 1182 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2746 6780 2774 6820
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 2455 6752 2774 6780
rect 2869 6783 2927 6789
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 2869 6743 2927 6749
rect 2884 6712 2912 6743
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3988 6780 4016 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 4617 6919 4675 6925
rect 4617 6885 4629 6919
rect 4663 6885 4675 6919
rect 4617 6879 4675 6885
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4246 6848 4252 6860
rect 4111 6820 4252 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 4632 6848 4660 6879
rect 8478 6848 8484 6860
rect 4580 6820 4660 6848
rect 4724 6820 8484 6848
rect 4580 6808 4586 6820
rect 3896 6752 4016 6780
rect 4157 6783 4215 6789
rect 3896 6712 3924 6752
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4724 6780 4752 6820
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 4203 6752 4752 6780
rect 4801 6783 4859 6789
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5718 6780 5724 6792
rect 5583 6752 5724 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 2884 6684 3924 6712
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4816 6712 4844 6743
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 18322 6780 18328 6792
rect 18283 6752 18328 6780
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 6454 6712 6460 6724
rect 4028 6684 4844 6712
rect 4908 6684 6460 6712
rect 4028 6672 4034 6684
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 1854 6644 1860 6656
rect 1811 6616 1860 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 4908 6644 4936 6684
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 3099 6616 4936 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 1762 6440 1768 6452
rect 1723 6412 1768 6440
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 2096 6412 3617 6440
rect 2096 6400 2102 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 3605 6403 3663 6409
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 4396 6412 4813 6440
rect 4396 6400 4402 6412
rect 4801 6409 4813 6412
rect 4847 6409 4859 6443
rect 4801 6403 4859 6409
rect 750 6332 756 6384
rect 808 6372 814 6384
rect 808 6344 2268 6372
rect 808 6332 814 6344
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 2240 6313 2268 6344
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 3016 6344 4384 6372
rect 3016 6332 3022 6344
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 900 6276 1593 6304
rect 900 6264 906 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 3510 6304 3516 6316
rect 2915 6276 3516 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 4356 6313 4384 6344
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4341 6307 4399 6313
rect 3743 6276 4200 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 658 6128 664 6180
rect 716 6168 722 6180
rect 4172 6177 4200 6276
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 4387 6276 5365 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 18322 6304 18328 6316
rect 18283 6276 18328 6304
rect 5353 6267 5411 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 2409 6171 2467 6177
rect 2409 6168 2421 6171
rect 716 6140 2421 6168
rect 716 6128 722 6140
rect 2409 6137 2421 6140
rect 2455 6137 2467 6171
rect 2409 6131 2467 6137
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6137 4215 6171
rect 4157 6131 4215 6137
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 1026 5856 1032 5908
rect 1084 5896 1090 5908
rect 2225 5899 2283 5905
rect 2225 5896 2237 5899
rect 1084 5868 2237 5896
rect 1084 5856 1090 5868
rect 2225 5865 2237 5868
rect 2271 5865 2283 5899
rect 2225 5859 2283 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3050 5896 3056 5908
rect 2915 5868 3056 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4617 5899 4675 5905
rect 4617 5896 4629 5899
rect 4028 5868 4629 5896
rect 4028 5856 4034 5868
rect 4617 5865 4629 5868
rect 4663 5865 4675 5899
rect 4617 5859 4675 5865
rect 1673 5831 1731 5837
rect 1673 5797 1685 5831
rect 1719 5828 1731 5831
rect 3602 5828 3608 5840
rect 1719 5800 3608 5828
rect 1719 5797 1731 5800
rect 1673 5791 1731 5797
rect 3602 5788 3608 5800
rect 3660 5788 3666 5840
rect 1210 5720 1216 5772
rect 1268 5760 1274 5772
rect 1268 5732 2452 5760
rect 1268 5720 1274 5732
rect 2424 5701 2452 5732
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 2409 5655 2467 5661
rect 1780 5624 1808 5655
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 4430 5624 4436 5636
rect 1780 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 1673 5355 1731 5361
rect 1673 5352 1685 5355
rect 1636 5324 1685 5352
rect 1636 5312 1642 5324
rect 1673 5321 1685 5324
rect 1719 5321 1731 5355
rect 1673 5315 1731 5321
rect 4522 5284 4528 5296
rect 1780 5256 4528 5284
rect 1780 5225 1808 5256
rect 4522 5244 4528 5256
rect 4580 5244 4586 5296
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2774 5216 2780 5228
rect 2271 5188 2780 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 2924 5188 2969 5216
rect 2924 5176 2930 5188
rect 18322 5080 18328 5092
rect 18283 5052 18328 5080
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 6086 4604 6092 4616
rect 1903 4576 6092 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19150 4604 19156 4616
rect 18371 4576 19156 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 18322 3924 18328 3936
rect 18283 3896 18328 3924
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 1578 3040 1584 3052
rect 1539 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 18322 2836 18328 2848
rect 18283 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 17678 2428 17684 2440
rect 17639 2400 17684 2428
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 9956 17688 10008 17740
rect 13544 17688 13596 17740
rect 8576 17620 8628 17672
rect 10508 17620 10560 17672
rect 6552 17552 6604 17604
rect 10600 17552 10652 17604
rect 5540 17484 5592 17536
rect 7104 17484 7156 17536
rect 9680 17484 9732 17536
rect 10692 17484 10744 17536
rect 13728 17484 13780 17536
rect 18788 17484 18840 17536
rect 19432 17484 19484 17536
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 9680 17280 9732 17332
rect 10600 17280 10652 17332
rect 11244 17280 11296 17332
rect 6552 17212 6604 17264
rect 10784 17212 10836 17264
rect 940 17144 992 17196
rect 5724 17144 5776 17196
rect 9128 17187 9180 17196
rect 1492 17076 1544 17128
rect 2964 17076 3016 17128
rect 5080 17008 5132 17060
rect 3516 16940 3568 16992
rect 3792 16940 3844 16992
rect 5172 16940 5224 16992
rect 5908 16940 5960 16992
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9312 17144 9364 17196
rect 9680 17144 9732 17196
rect 11060 17144 11112 17196
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 15200 17187 15252 17196
rect 15200 17153 15234 17187
rect 15234 17153 15252 17187
rect 15200 17144 15252 17153
rect 17960 17144 18012 17196
rect 10324 17076 10376 17128
rect 10508 17076 10560 17128
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 16948 17119 17000 17128
rect 16948 17085 16957 17119
rect 16957 17085 16991 17119
rect 16991 17085 17000 17119
rect 16948 17076 17000 17085
rect 6000 16940 6052 16949
rect 6828 16940 6880 16992
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 10416 17008 10468 17060
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 16304 16983 16356 16992
rect 16304 16949 16313 16983
rect 16313 16949 16347 16983
rect 16347 16949 16356 16983
rect 16304 16940 16356 16949
rect 17132 16940 17184 16992
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 11152 16736 11204 16788
rect 11612 16736 11664 16788
rect 12348 16779 12400 16788
rect 3516 16668 3568 16720
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 12624 16736 12676 16788
rect 2964 16643 3016 16652
rect 1676 16532 1728 16584
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 3884 16532 3936 16584
rect 3332 16464 3384 16516
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 4252 16507 4304 16516
rect 4252 16473 4261 16507
rect 4261 16473 4295 16507
rect 4295 16473 4304 16507
rect 4252 16464 4304 16473
rect 6644 16600 6696 16652
rect 13084 16668 13136 16720
rect 15844 16736 15896 16788
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 6828 16532 6880 16584
rect 6184 16464 6236 16516
rect 6552 16507 6604 16516
rect 6552 16473 6561 16507
rect 6561 16473 6595 16507
rect 6595 16473 6604 16507
rect 6552 16464 6604 16473
rect 7288 16532 7340 16584
rect 8944 16532 8996 16584
rect 4436 16396 4488 16448
rect 4896 16396 4948 16448
rect 4988 16439 5040 16448
rect 4988 16405 4997 16439
rect 4997 16405 5031 16439
rect 5031 16405 5040 16439
rect 4988 16396 5040 16405
rect 7288 16396 7340 16448
rect 8668 16464 8720 16516
rect 10232 16507 10284 16516
rect 10232 16473 10250 16507
rect 10250 16473 10284 16507
rect 10232 16464 10284 16473
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 10692 16532 10744 16584
rect 11428 16464 11480 16516
rect 11704 16532 11756 16584
rect 14280 16532 14332 16584
rect 15016 16532 15068 16584
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 16212 16532 16264 16584
rect 17132 16532 17184 16584
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17776 16575 17828 16584
rect 17408 16532 17460 16541
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 12348 16464 12400 16516
rect 13268 16507 13320 16516
rect 13268 16473 13277 16507
rect 13277 16473 13311 16507
rect 13311 16473 13320 16507
rect 13268 16464 13320 16473
rect 13912 16464 13964 16516
rect 15292 16464 15344 16516
rect 16120 16464 16172 16516
rect 7656 16396 7708 16448
rect 8300 16396 8352 16448
rect 8392 16396 8444 16448
rect 9588 16396 9640 16448
rect 10968 16396 11020 16448
rect 11796 16396 11848 16448
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 3884 16192 3936 16244
rect 4528 16192 4580 16244
rect 6000 16192 6052 16244
rect 6920 16192 6972 16244
rect 10968 16192 11020 16244
rect 11152 16192 11204 16244
rect 3332 16124 3384 16176
rect 1676 16056 1728 16108
rect 2228 16056 2280 16108
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 3884 16056 3936 16108
rect 4344 16124 4396 16176
rect 6552 16124 6604 16176
rect 7288 16124 7340 16176
rect 7656 16124 7708 16176
rect 8024 16167 8076 16176
rect 8024 16133 8029 16167
rect 8029 16133 8063 16167
rect 8063 16133 8076 16167
rect 8024 16124 8076 16133
rect 8300 16124 8352 16176
rect 4712 16056 4764 16108
rect 7196 16056 7248 16108
rect 8668 16056 8720 16108
rect 8852 16056 8904 16108
rect 9036 16099 9088 16108
rect 9036 16065 9070 16099
rect 9070 16065 9088 16099
rect 9036 16056 9088 16065
rect 9588 16056 9640 16108
rect 10784 16099 10836 16108
rect 4068 15988 4120 16040
rect 5724 15988 5776 16040
rect 8300 15988 8352 16040
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 12256 16124 12308 16176
rect 11520 16056 11572 16108
rect 13452 16124 13504 16176
rect 14556 16192 14608 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 14372 16124 14424 16176
rect 15384 16124 15436 16176
rect 17408 16124 17460 16176
rect 3608 15920 3660 15972
rect 4252 15920 4304 15972
rect 4436 15963 4488 15972
rect 4436 15929 4445 15963
rect 4445 15929 4479 15963
rect 4479 15929 4488 15963
rect 4436 15920 4488 15929
rect 3056 15852 3108 15904
rect 3700 15852 3752 15904
rect 3976 15852 4028 15904
rect 4988 15920 5040 15972
rect 5172 15920 5224 15972
rect 6092 15920 6144 15972
rect 6828 15920 6880 15972
rect 11888 15988 11940 16040
rect 12256 15988 12308 16040
rect 12900 15988 12952 16040
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 7840 15852 7892 15904
rect 11796 15963 11848 15972
rect 11796 15929 11805 15963
rect 11805 15929 11839 15963
rect 11839 15929 11848 15963
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 11796 15920 11848 15929
rect 9496 15852 9548 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 12440 15852 12492 15904
rect 13176 15920 13228 15972
rect 14096 15988 14148 16040
rect 16304 16056 16356 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 14924 16031 14976 16040
rect 14924 15997 14933 16031
rect 14933 15997 14967 16031
rect 14967 15997 14976 16031
rect 14924 15988 14976 15997
rect 15936 15988 15988 16040
rect 14740 15852 14792 15904
rect 14924 15852 14976 15904
rect 16856 15852 16908 15904
rect 18052 15852 18104 15904
rect 19248 15852 19300 15904
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 1492 15648 1544 15700
rect 664 15580 716 15632
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 3056 15512 3108 15564
rect 3700 15512 3752 15564
rect 4896 15648 4948 15700
rect 5080 15444 5132 15496
rect 7104 15648 7156 15700
rect 7564 15648 7616 15700
rect 7288 15580 7340 15632
rect 7840 15580 7892 15632
rect 6460 15512 6512 15564
rect 9128 15648 9180 15700
rect 9220 15648 9272 15700
rect 8024 15580 8076 15632
rect 8392 15580 8444 15632
rect 8760 15580 8812 15632
rect 10508 15580 10560 15632
rect 12716 15648 12768 15700
rect 13268 15648 13320 15700
rect 14832 15648 14884 15700
rect 15016 15691 15068 15700
rect 15016 15657 15025 15691
rect 15025 15657 15059 15691
rect 15059 15657 15068 15691
rect 15016 15648 15068 15657
rect 6736 15444 6788 15496
rect 1952 15308 2004 15360
rect 3056 15376 3108 15428
rect 3884 15376 3936 15428
rect 6920 15376 6972 15428
rect 7748 15444 7800 15496
rect 8944 15512 8996 15564
rect 12164 15580 12216 15632
rect 13544 15623 13596 15632
rect 13544 15589 13553 15623
rect 13553 15589 13587 15623
rect 13587 15589 13596 15623
rect 13544 15580 13596 15589
rect 14004 15580 14056 15632
rect 15384 15648 15436 15700
rect 15936 15648 15988 15700
rect 17868 15648 17920 15700
rect 8116 15376 8168 15428
rect 9680 15444 9732 15496
rect 8760 15376 8812 15428
rect 10692 15444 10744 15496
rect 10876 15376 10928 15428
rect 5172 15308 5224 15360
rect 5816 15308 5868 15360
rect 6644 15308 6696 15360
rect 7196 15308 7248 15360
rect 8944 15308 8996 15360
rect 9312 15308 9364 15360
rect 10692 15308 10744 15360
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 11244 15512 11296 15564
rect 12072 15512 12124 15564
rect 12716 15512 12768 15564
rect 12992 15512 13044 15564
rect 13268 15444 13320 15496
rect 11796 15376 11848 15428
rect 12440 15376 12492 15428
rect 12992 15376 13044 15428
rect 14556 15512 14608 15564
rect 15292 15580 15344 15632
rect 18052 15580 18104 15632
rect 15016 15444 15068 15496
rect 15936 15487 15988 15496
rect 14096 15376 14148 15428
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16212 15444 16264 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 16856 15376 16908 15428
rect 17776 15444 17828 15496
rect 17224 15419 17276 15428
rect 17224 15385 17258 15419
rect 17258 15385 17276 15419
rect 17224 15376 17276 15385
rect 12532 15308 12584 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 13636 15308 13688 15360
rect 13728 15308 13780 15360
rect 15752 15308 15804 15360
rect 18420 15376 18472 15428
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 3608 15104 3660 15156
rect 4896 15104 4948 15156
rect 5080 15147 5132 15156
rect 5080 15113 5089 15147
rect 5089 15113 5123 15147
rect 5123 15113 5132 15147
rect 5080 15104 5132 15113
rect 1676 14968 1728 15020
rect 2320 14968 2372 15020
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3976 15011 4028 15020
rect 3792 14968 3844 14977
rect 3976 14977 3984 15011
rect 3984 14977 4018 15011
rect 4018 14977 4028 15011
rect 3976 14968 4028 14977
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4528 15011 4580 15020
rect 4068 14968 4120 14977
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4988 15036 5040 15088
rect 5540 15079 5592 15088
rect 5540 15045 5549 15079
rect 5549 15045 5583 15079
rect 5583 15045 5592 15079
rect 5540 15036 5592 15045
rect 6000 15036 6052 15088
rect 8760 15104 8812 15156
rect 9404 15104 9456 15156
rect 7288 15036 7340 15088
rect 8116 15036 8168 15088
rect 8300 15036 8352 15088
rect 9864 15036 9916 15088
rect 5356 14968 5408 15020
rect 5080 14900 5132 14952
rect 5448 14900 5500 14952
rect 9680 14968 9732 15020
rect 10784 15104 10836 15156
rect 10968 15036 11020 15088
rect 12808 15104 12860 15156
rect 14556 15104 14608 15156
rect 15936 15104 15988 15156
rect 17408 15104 17460 15156
rect 12072 15079 12124 15088
rect 5816 14832 5868 14884
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 4896 14764 4948 14816
rect 8024 14900 8076 14952
rect 8116 14900 8168 14952
rect 9588 14900 9640 14952
rect 11244 14968 11296 15020
rect 11704 14900 11756 14952
rect 7564 14832 7616 14884
rect 6736 14764 6788 14816
rect 7472 14764 7524 14816
rect 10508 14832 10560 14884
rect 10692 14832 10744 14884
rect 12072 15045 12081 15079
rect 12081 15045 12115 15079
rect 12115 15045 12124 15079
rect 12072 15036 12124 15045
rect 13176 15036 13228 15088
rect 11980 14968 12032 15020
rect 14346 15079 14398 15088
rect 14346 15045 14355 15079
rect 14355 15045 14389 15079
rect 14389 15045 14398 15079
rect 14346 15036 14398 15045
rect 16304 15036 16356 15088
rect 17776 15036 17828 15088
rect 15568 14900 15620 14952
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 16212 14968 16264 15020
rect 18052 14968 18104 15020
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 14556 14832 14608 14884
rect 8576 14807 8628 14816
rect 8576 14773 8585 14807
rect 8585 14773 8619 14807
rect 8619 14773 8628 14807
rect 8576 14764 8628 14773
rect 8852 14764 8904 14816
rect 11152 14764 11204 14816
rect 11796 14764 11848 14816
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 14648 14764 14700 14816
rect 15384 14764 15436 14816
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 16396 14764 16448 14816
rect 18144 14764 18196 14816
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 756 14560 808 14612
rect 3884 14560 3936 14612
rect 4436 14560 4488 14612
rect 5172 14560 5224 14612
rect 7288 14560 7340 14612
rect 8392 14603 8444 14612
rect 4620 14492 4672 14544
rect 5448 14492 5500 14544
rect 5908 14492 5960 14544
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 10324 14560 10376 14612
rect 10508 14560 10560 14612
rect 11244 14560 11296 14612
rect 12440 14603 12492 14612
rect 1676 14356 1728 14408
rect 4988 14424 5040 14476
rect 5540 14424 5592 14476
rect 4344 14356 4396 14408
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 3424 14288 3476 14340
rect 3056 14220 3108 14272
rect 3976 14220 4028 14272
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4528 14220 4580 14272
rect 5264 14288 5316 14340
rect 5448 14288 5500 14340
rect 5816 14220 5868 14272
rect 6092 14220 6144 14272
rect 6920 14399 6972 14408
rect 6920 14365 6929 14399
rect 6929 14365 6963 14399
rect 6963 14365 6972 14399
rect 7564 14492 7616 14544
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13820 14560 13872 14612
rect 15016 14560 15068 14612
rect 15200 14560 15252 14612
rect 15384 14560 15436 14612
rect 8208 14424 8260 14476
rect 9864 14424 9916 14476
rect 10324 14424 10376 14476
rect 13084 14492 13136 14544
rect 13176 14492 13228 14544
rect 16948 14560 17000 14612
rect 17500 14560 17552 14612
rect 17132 14492 17184 14544
rect 13452 14424 13504 14476
rect 15844 14424 15896 14476
rect 6920 14356 6972 14365
rect 8852 14356 8904 14408
rect 9128 14356 9180 14408
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 10600 14356 10652 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 15384 14356 15436 14408
rect 15568 14356 15620 14408
rect 7196 14288 7248 14340
rect 7840 14288 7892 14340
rect 9588 14288 9640 14340
rect 11704 14331 11756 14340
rect 11704 14297 11722 14331
rect 11722 14297 11756 14331
rect 11704 14288 11756 14297
rect 12900 14288 12952 14340
rect 14372 14288 14424 14340
rect 15200 14288 15252 14340
rect 16304 14356 16356 14408
rect 18144 14424 18196 14476
rect 18236 14399 18288 14408
rect 18236 14365 18244 14399
rect 18244 14365 18278 14399
rect 18278 14365 18288 14399
rect 18236 14356 18288 14365
rect 8852 14220 8904 14272
rect 9404 14220 9456 14272
rect 11244 14220 11296 14272
rect 11336 14220 11388 14272
rect 12532 14220 12584 14272
rect 16212 14220 16264 14272
rect 16764 14220 16816 14272
rect 17040 14220 17092 14272
rect 18144 14288 18196 14340
rect 18052 14220 18104 14272
rect 18328 14220 18380 14272
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 3424 14016 3476 14068
rect 3884 14059 3936 14068
rect 3884 14025 3893 14059
rect 3893 14025 3927 14059
rect 3927 14025 3936 14059
rect 3884 14016 3936 14025
rect 7840 14016 7892 14068
rect 9128 14016 9180 14068
rect 9680 14016 9732 14068
rect 9956 14016 10008 14068
rect 10140 14016 10192 14068
rect 11336 14016 11388 14068
rect 11704 14059 11756 14068
rect 11704 14025 11713 14059
rect 11713 14025 11747 14059
rect 11747 14025 11756 14059
rect 11704 14016 11756 14025
rect 13912 14016 13964 14068
rect 14280 14016 14332 14068
rect 14648 14016 14700 14068
rect 16580 14016 16632 14068
rect 1952 13948 2004 14000
rect 4160 13948 4212 14000
rect 5264 13948 5316 14000
rect 1492 13880 1544 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 5080 13880 5132 13932
rect 5356 13880 5408 13932
rect 2596 13744 2648 13796
rect 3792 13744 3844 13796
rect 4160 13812 4212 13864
rect 5632 13812 5684 13864
rect 5080 13744 5132 13796
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 4528 13676 4580 13685
rect 6920 13948 6972 14000
rect 8484 13948 8536 14000
rect 8576 13948 8628 14000
rect 8852 13948 8904 14000
rect 6644 13880 6696 13932
rect 8208 13880 8260 13932
rect 9128 13880 9180 13932
rect 11520 13948 11572 14000
rect 15200 13948 15252 14000
rect 11244 13880 11296 13932
rect 13728 13880 13780 13932
rect 14188 13880 14240 13932
rect 16212 13948 16264 14000
rect 16488 13948 16540 14000
rect 16948 13948 17000 14000
rect 17408 13948 17460 14000
rect 18144 14016 18196 14068
rect 15936 13880 15988 13932
rect 6460 13812 6512 13864
rect 7840 13812 7892 13864
rect 8116 13812 8168 13864
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 9496 13744 9548 13796
rect 11796 13812 11848 13864
rect 9772 13744 9824 13796
rect 10416 13744 10468 13796
rect 14372 13812 14424 13864
rect 15476 13787 15528 13796
rect 15476 13753 15485 13787
rect 15485 13753 15519 13787
rect 15519 13753 15528 13787
rect 15476 13744 15528 13753
rect 8208 13676 8260 13728
rect 8484 13676 8536 13728
rect 10140 13676 10192 13728
rect 12624 13676 12676 13728
rect 14556 13676 14608 13728
rect 16304 13812 16356 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 16764 13744 16816 13796
rect 17408 13812 17460 13864
rect 18512 13744 18564 13796
rect 16672 13676 16724 13728
rect 18236 13676 18288 13728
rect 18696 13676 18748 13728
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 4160 13515 4212 13524
rect 2596 13404 2648 13456
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 5816 13515 5868 13524
rect 5816 13481 5825 13515
rect 5825 13481 5859 13515
rect 5859 13481 5868 13515
rect 5816 13472 5868 13481
rect 6000 13515 6052 13524
rect 6000 13481 6009 13515
rect 6009 13481 6043 13515
rect 6043 13481 6052 13515
rect 6644 13515 6696 13524
rect 6000 13472 6052 13481
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 6828 13472 6880 13524
rect 1952 13336 2004 13388
rect 3516 13336 3568 13388
rect 5632 13336 5684 13388
rect 1216 13200 1268 13252
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 3976 13243 4028 13252
rect 3976 13209 3985 13243
rect 3985 13209 4019 13243
rect 4019 13209 4028 13243
rect 3976 13200 4028 13209
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 4620 13132 4672 13184
rect 4896 13200 4948 13252
rect 6184 13200 6236 13252
rect 7472 13472 7524 13524
rect 7656 13472 7708 13524
rect 11520 13472 11572 13524
rect 11888 13472 11940 13524
rect 16948 13472 17000 13524
rect 17316 13472 17368 13524
rect 18696 13472 18748 13524
rect 7748 13404 7800 13456
rect 9496 13404 9548 13456
rect 7104 13268 7156 13320
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 7380 13200 7432 13252
rect 8208 13336 8260 13388
rect 9404 13336 9456 13388
rect 9864 13336 9916 13388
rect 10968 13404 11020 13456
rect 18144 13447 18196 13456
rect 13268 13336 13320 13388
rect 13544 13336 13596 13388
rect 14740 13336 14792 13388
rect 8576 13268 8628 13320
rect 9312 13268 9364 13320
rect 10416 13268 10468 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 5356 13132 5408 13184
rect 6000 13132 6052 13184
rect 7472 13132 7524 13184
rect 8484 13200 8536 13252
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 9956 13132 10008 13184
rect 11520 13268 11572 13320
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 12900 13268 12952 13277
rect 15108 13268 15160 13320
rect 15292 13268 15344 13320
rect 17132 13336 17184 13388
rect 15752 13268 15804 13320
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 16396 13268 16448 13320
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 18144 13413 18153 13447
rect 18153 13413 18187 13447
rect 18187 13413 18196 13447
rect 18144 13404 18196 13413
rect 17040 13268 17092 13277
rect 17132 13200 17184 13252
rect 13360 13132 13412 13184
rect 15200 13132 15252 13184
rect 16212 13132 16264 13184
rect 18512 13132 18564 13184
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 1308 12928 1360 12980
rect 4804 12928 4856 12980
rect 5080 12928 5132 12980
rect 7564 12928 7616 12980
rect 2688 12860 2740 12912
rect 4252 12860 4304 12912
rect 4528 12903 4580 12912
rect 4528 12869 4537 12903
rect 4537 12869 4571 12903
rect 4571 12869 4580 12903
rect 4528 12860 4580 12869
rect 6460 12860 6512 12912
rect 8760 12928 8812 12980
rect 10232 12928 10284 12980
rect 10876 12928 10928 12980
rect 11612 12928 11664 12980
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 3792 12792 3844 12844
rect 8852 12792 8904 12844
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 4804 12724 4856 12776
rect 3700 12656 3752 12708
rect 4344 12588 4396 12640
rect 4712 12656 4764 12708
rect 6092 12724 6144 12776
rect 7656 12724 7708 12776
rect 9496 12792 9548 12844
rect 9588 12792 9640 12844
rect 10784 12792 10836 12844
rect 10968 12792 11020 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 13452 12928 13504 12980
rect 17868 12971 17920 12980
rect 17868 12937 17877 12971
rect 17877 12937 17911 12971
rect 17911 12937 17920 12971
rect 17868 12928 17920 12937
rect 18144 12928 18196 12980
rect 18328 12928 18380 12980
rect 13912 12860 13964 12912
rect 14740 12860 14792 12912
rect 17408 12903 17460 12912
rect 17408 12869 17417 12903
rect 17417 12869 17451 12903
rect 17451 12869 17460 12903
rect 17408 12860 17460 12869
rect 9404 12724 9456 12776
rect 11244 12724 11296 12776
rect 13820 12792 13872 12844
rect 14648 12792 14700 12844
rect 14924 12792 14976 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 16396 12792 16448 12844
rect 17776 12792 17828 12844
rect 15200 12724 15252 12776
rect 16212 12724 16264 12776
rect 5632 12656 5684 12708
rect 6460 12656 6512 12708
rect 7564 12656 7616 12708
rect 11796 12656 11848 12708
rect 15476 12699 15528 12708
rect 15476 12665 15485 12699
rect 15485 12665 15519 12699
rect 15519 12665 15528 12699
rect 15476 12656 15528 12665
rect 16304 12699 16356 12708
rect 16304 12665 16313 12699
rect 16313 12665 16347 12699
rect 16347 12665 16356 12699
rect 16304 12656 16356 12665
rect 6920 12588 6972 12640
rect 7472 12588 7524 12640
rect 9404 12588 9456 12640
rect 10140 12588 10192 12640
rect 14004 12588 14056 12640
rect 14832 12588 14884 12640
rect 16856 12588 16908 12640
rect 17960 12656 18012 12708
rect 18328 12656 18380 12708
rect 18512 12656 18564 12708
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 2872 12384 2924 12436
rect 4620 12384 4672 12436
rect 6552 12427 6604 12436
rect 6552 12393 6561 12427
rect 6561 12393 6595 12427
rect 6595 12393 6604 12427
rect 6552 12384 6604 12393
rect 6828 12384 6880 12436
rect 9036 12384 9088 12436
rect 9772 12384 9824 12436
rect 11060 12384 11112 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 15016 12384 15068 12436
rect 940 12248 992 12300
rect 1308 12248 1360 12300
rect 1492 12248 1544 12300
rect 3792 12248 3844 12300
rect 1308 12112 1360 12164
rect 1768 12044 1820 12096
rect 3700 12112 3752 12164
rect 4068 12112 4120 12164
rect 6644 12316 6696 12368
rect 6736 12316 6788 12368
rect 4988 12155 5040 12164
rect 4988 12121 5015 12155
rect 5015 12121 5040 12155
rect 2964 12087 3016 12096
rect 2964 12053 2973 12087
rect 2973 12053 3007 12087
rect 3007 12053 3016 12087
rect 2964 12044 3016 12053
rect 3424 12044 3476 12096
rect 4988 12112 5040 12121
rect 5080 12112 5132 12164
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 6000 12180 6052 12232
rect 6184 12112 6236 12164
rect 6368 12112 6420 12164
rect 6828 12180 6880 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 8300 12180 8352 12232
rect 8484 12248 8536 12300
rect 9128 12316 9180 12368
rect 10876 12316 10928 12368
rect 16396 12316 16448 12368
rect 16948 12384 17000 12436
rect 17500 12384 17552 12436
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 19248 12316 19300 12368
rect 10416 12248 10468 12300
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 8944 12180 8996 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 12808 12248 12860 12300
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11244 12180 11296 12232
rect 15844 12248 15896 12300
rect 16028 12291 16080 12300
rect 16028 12257 16037 12291
rect 16037 12257 16071 12291
rect 16071 12257 16080 12291
rect 16028 12248 16080 12257
rect 17408 12248 17460 12300
rect 7472 12112 7524 12164
rect 7656 12044 7708 12096
rect 12992 12112 13044 12164
rect 15016 12112 15068 12164
rect 15292 12180 15344 12232
rect 16304 12180 16356 12232
rect 17040 12112 17092 12164
rect 17316 12155 17368 12164
rect 17316 12121 17325 12155
rect 17325 12121 17359 12155
rect 17359 12121 17368 12155
rect 17316 12112 17368 12121
rect 17408 12112 17460 12164
rect 10692 12044 10744 12096
rect 16396 12044 16448 12096
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 2872 11840 2924 11892
rect 4436 11840 4488 11892
rect 4528 11840 4580 11892
rect 6552 11840 6604 11892
rect 7748 11840 7800 11892
rect 9404 11840 9456 11892
rect 9680 11840 9732 11892
rect 10232 11840 10284 11892
rect 10416 11840 10468 11892
rect 10876 11883 10928 11892
rect 1492 11704 1544 11756
rect 2136 11704 2188 11756
rect 3516 11772 3568 11824
rect 4988 11772 5040 11824
rect 3608 11636 3660 11688
rect 4712 11704 4764 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5264 11704 5316 11756
rect 5724 11815 5776 11824
rect 5724 11781 5733 11815
rect 5733 11781 5767 11815
rect 5767 11781 5776 11815
rect 5724 11772 5776 11781
rect 7656 11772 7708 11824
rect 9496 11772 9548 11824
rect 6460 11704 6512 11756
rect 7012 11704 7064 11756
rect 7932 11704 7984 11756
rect 8668 11704 8720 11756
rect 10600 11772 10652 11824
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 14096 11840 14148 11892
rect 15476 11840 15528 11892
rect 17408 11840 17460 11892
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 10876 11747 10928 11756
rect 3884 11636 3936 11688
rect 848 11568 900 11620
rect 1124 11568 1176 11620
rect 3424 11500 3476 11552
rect 4068 11500 4120 11552
rect 4252 11500 4304 11552
rect 5080 11636 5132 11688
rect 7288 11636 7340 11688
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 15016 11772 15068 11824
rect 19432 11840 19484 11892
rect 18328 11815 18380 11824
rect 18328 11781 18337 11815
rect 18337 11781 18371 11815
rect 18371 11781 18380 11815
rect 18328 11772 18380 11781
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 14648 11704 14700 11756
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 15292 11704 15344 11756
rect 5356 11611 5408 11620
rect 5356 11577 5365 11611
rect 5365 11577 5399 11611
rect 5399 11577 5408 11611
rect 5356 11568 5408 11577
rect 7932 11568 7984 11620
rect 14740 11636 14792 11688
rect 15936 11704 15988 11756
rect 17960 11704 18012 11756
rect 18052 11636 18104 11688
rect 9404 11568 9456 11620
rect 11428 11568 11480 11620
rect 17500 11611 17552 11620
rect 17500 11577 17509 11611
rect 17509 11577 17543 11611
rect 17543 11577 17552 11611
rect 17500 11568 17552 11577
rect 5080 11500 5132 11552
rect 5724 11500 5776 11552
rect 6276 11500 6328 11552
rect 10876 11500 10928 11552
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 1124 11296 1176 11348
rect 5264 11296 5316 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 7472 11296 7524 11348
rect 9680 11296 9732 11348
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14188 11296 14240 11348
rect 16120 11296 16172 11348
rect 17132 11296 17184 11348
rect 17316 11296 17368 11348
rect 3516 11228 3568 11280
rect 4344 11228 4396 11280
rect 5172 11228 5224 11280
rect 5356 11228 5408 11280
rect 8116 11228 8168 11280
rect 11060 11271 11112 11280
rect 1492 11160 1544 11212
rect 2872 11160 2924 11212
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 5080 11092 5132 11144
rect 5172 11092 5224 11144
rect 5908 11160 5960 11212
rect 6184 11160 6236 11212
rect 1860 11067 1912 11076
rect 1860 11033 1894 11067
rect 1894 11033 1912 11067
rect 1860 11024 1912 11033
rect 2504 11024 2556 11076
rect 5908 11067 5960 11076
rect 5908 11033 5917 11067
rect 5917 11033 5951 11067
rect 5951 11033 5960 11067
rect 5908 11024 5960 11033
rect 6276 11092 6328 11144
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 8116 11135 8168 11144
rect 6736 11024 6788 11076
rect 2688 10956 2740 11008
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 5172 10956 5224 11008
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 11060 11237 11069 11271
rect 11069 11237 11103 11271
rect 11103 11237 11112 11271
rect 11060 11228 11112 11237
rect 14464 11271 14516 11280
rect 14464 11237 14473 11271
rect 14473 11237 14507 11271
rect 14507 11237 14516 11271
rect 14464 11228 14516 11237
rect 14924 11228 14976 11280
rect 17684 11228 17736 11280
rect 9496 11160 9548 11212
rect 16396 11135 16448 11144
rect 16396 11101 16405 11135
rect 16405 11101 16439 11135
rect 16439 11101 16448 11135
rect 16396 11092 16448 11101
rect 17132 11160 17184 11212
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17868 11092 17920 11144
rect 18512 11092 18564 11144
rect 17408 11024 17460 11076
rect 13268 10956 13320 11008
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 2228 10752 2280 10804
rect 6920 10795 6972 10804
rect 2964 10684 3016 10736
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 10324 10752 10376 10804
rect 15108 10752 15160 10804
rect 17224 10752 17276 10804
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 1584 10480 1636 10532
rect 2688 10616 2740 10668
rect 2228 10412 2280 10464
rect 3792 10616 3844 10668
rect 3976 10616 4028 10668
rect 4528 10616 4580 10668
rect 5540 10616 5592 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7380 10659 7432 10668
rect 5356 10548 5408 10600
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 9220 10616 9272 10668
rect 9588 10616 9640 10668
rect 15752 10616 15804 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 18420 10684 18472 10736
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 7288 10548 7340 10600
rect 8116 10548 8168 10600
rect 18604 10548 18656 10600
rect 5908 10480 5960 10532
rect 18236 10480 18288 10532
rect 2412 10412 2464 10464
rect 2596 10412 2648 10464
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 2780 10208 2832 10260
rect 4528 10208 4580 10260
rect 5080 10208 5132 10260
rect 5264 10208 5316 10260
rect 5540 10208 5592 10260
rect 6552 10208 6604 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 8024 10208 8076 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9312 10208 9364 10260
rect 15384 10208 15436 10260
rect 1492 10072 1544 10124
rect 2412 10004 2464 10056
rect 2228 9936 2280 9988
rect 1952 9868 2004 9920
rect 2964 10072 3016 10124
rect 3056 10072 3108 10124
rect 5080 10072 5132 10124
rect 4252 10047 4304 10056
rect 3056 9936 3108 9988
rect 3424 9868 3476 9920
rect 3792 9868 3844 9920
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 4712 10004 4764 10056
rect 4988 10004 5040 10056
rect 4160 9936 4212 9988
rect 5448 9936 5500 9988
rect 6644 10004 6696 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 9680 10004 9732 10056
rect 16212 10208 16264 10260
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 15568 10140 15620 10192
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 10508 9936 10560 9988
rect 4436 9868 4488 9920
rect 4620 9868 4672 9920
rect 5264 9868 5316 9920
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 2872 9664 2924 9716
rect 2412 9596 2464 9648
rect 2596 9596 2648 9648
rect 3516 9528 3568 9580
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3792 9571 3844 9580
rect 3608 9528 3660 9537
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 2780 9460 2832 9512
rect 4160 9596 4212 9648
rect 4620 9596 4672 9648
rect 4896 9639 4948 9648
rect 4896 9605 4905 9639
rect 4905 9605 4939 9639
rect 4939 9605 4948 9639
rect 4896 9596 4948 9605
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 5908 9664 5960 9716
rect 7564 9664 7616 9716
rect 9680 9596 9732 9648
rect 17684 9664 17736 9716
rect 4068 9528 4120 9580
rect 5356 9571 5408 9580
rect 4160 9460 4212 9512
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 3884 9392 3936 9444
rect 4344 9392 4396 9444
rect 4620 9435 4672 9444
rect 4620 9401 4629 9435
rect 4629 9401 4663 9435
rect 4663 9401 4672 9435
rect 4620 9392 4672 9401
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 5448 9528 5500 9580
rect 4988 9460 5040 9512
rect 8208 9528 8260 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 17960 9596 18012 9648
rect 19064 9596 19116 9648
rect 15200 9460 15252 9512
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 14648 9392 14700 9444
rect 19156 9460 19208 9512
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 2320 9120 2372 9172
rect 4988 9120 5040 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 7012 9120 7064 9172
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 8668 9120 8720 9172
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 3700 9052 3752 9104
rect 4528 9052 4580 9104
rect 8024 9052 8076 9104
rect 17868 9052 17920 9104
rect 3056 8984 3108 9036
rect 1952 8848 2004 8900
rect 2596 8848 2648 8900
rect 2872 8848 2924 8900
rect 2412 8780 2464 8832
rect 5448 8984 5500 9036
rect 17960 8984 18012 9036
rect 4160 8916 4212 8968
rect 4804 8916 4856 8968
rect 5356 8916 5408 8968
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 7104 8916 7156 8968
rect 3424 8848 3476 8900
rect 4252 8848 4304 8900
rect 4620 8848 4672 8900
rect 5908 8848 5960 8900
rect 3884 8780 3936 8832
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 2320 8576 2372 8628
rect 2412 8576 2464 8628
rect 3332 8576 3384 8628
rect 1676 8508 1728 8560
rect 2688 8508 2740 8560
rect 2596 8440 2648 8492
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 2688 8372 2740 8424
rect 3424 8440 3476 8492
rect 7932 8576 7984 8628
rect 17592 8576 17644 8628
rect 4160 8440 4212 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 5724 8440 5776 8492
rect 7196 8483 7248 8492
rect 3700 8372 3752 8424
rect 4068 8372 4120 8424
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 19156 8440 19208 8492
rect 2320 8236 2372 8288
rect 3424 8236 3476 8288
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 4436 8304 4488 8356
rect 4620 8236 4672 8288
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 2688 8032 2740 8084
rect 3976 8075 4028 8084
rect 3976 8041 3985 8075
rect 3985 8041 4019 8075
rect 4019 8041 4028 8075
rect 3976 8032 4028 8041
rect 4712 8075 4764 8084
rect 4712 8041 4721 8075
rect 4721 8041 4755 8075
rect 4755 8041 4764 8075
rect 4712 8032 4764 8041
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 9588 8032 9640 8084
rect 1584 7828 1636 7880
rect 3792 7964 3844 8016
rect 6552 7964 6604 8016
rect 1952 7828 2004 7880
rect 2320 7828 2372 7880
rect 3056 7828 3108 7880
rect 5632 7896 5684 7948
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 7104 7828 7156 7880
rect 2780 7803 2832 7812
rect 2780 7769 2807 7803
rect 2807 7769 2832 7803
rect 2780 7760 2832 7769
rect 572 7692 624 7744
rect 2320 7692 2372 7744
rect 2412 7692 2464 7744
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 2136 7488 2188 7540
rect 2872 7488 2924 7540
rect 1676 7420 1728 7472
rect 5080 7488 5132 7540
rect 5816 7488 5868 7540
rect 6184 7488 6236 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 6000 7420 6052 7472
rect 940 7216 992 7268
rect 5816 7395 5868 7404
rect 1308 7148 1360 7200
rect 3148 7284 3200 7336
rect 4068 7284 4120 7336
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 6368 7284 6420 7336
rect 2320 7216 2372 7268
rect 5908 7216 5960 7268
rect 6276 7148 6328 7200
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 5816 6944 5868 6996
rect 1124 6740 1176 6792
rect 3884 6808 3936 6860
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 4160 6876 4212 6928
rect 4252 6808 4304 6860
rect 4528 6808 4580 6860
rect 8484 6808 8536 6860
rect 3976 6672 4028 6724
rect 5724 6740 5776 6792
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 1860 6604 1912 6656
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 6460 6672 6512 6724
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2044 6400 2096 6452
rect 4344 6400 4396 6452
rect 756 6332 808 6384
rect 848 6264 900 6316
rect 2964 6332 3016 6384
rect 3516 6264 3568 6316
rect 664 6128 716 6180
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 1032 5856 1084 5908
rect 3056 5856 3108 5908
rect 3976 5856 4028 5908
rect 3608 5788 3660 5840
rect 1216 5720 1268 5772
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 4436 5584 4488 5636
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 1584 5312 1636 5364
rect 4528 5244 4580 5296
rect 2780 5176 2832 5228
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 18328 5083 18380 5092
rect 18328 5049 18337 5083
rect 18337 5049 18371 5083
rect 18371 5049 18380 5083
rect 18328 5040 18380 5049
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 6092 4564 6144 4616
rect 19156 4564 19208 4616
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 386 19200 442 20000
rect 584 19230 1072 19258
rect 400 18601 428 19200
rect 386 18592 442 18601
rect 386 18527 442 18536
rect 584 7750 612 19230
rect 1044 19122 1072 19230
rect 1122 19200 1178 20000
rect 1858 19200 1914 20000
rect 2594 19200 2650 20000
rect 3330 19200 3386 20000
rect 3436 19230 3740 19258
rect 1136 19122 1164 19200
rect 1044 19094 1164 19122
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 16574 980 17138
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 952 16546 1072 16574
rect 664 15632 716 15638
rect 664 15574 716 15580
rect 572 7744 624 7750
rect 572 7686 624 7692
rect 676 6186 704 15574
rect 756 14612 808 14618
rect 756 14554 808 14560
rect 768 6390 796 14554
rect 940 12300 992 12306
rect 940 12242 992 12248
rect 848 11620 900 11626
rect 848 11562 900 11568
rect 756 6384 808 6390
rect 756 6326 808 6332
rect 860 6322 888 11562
rect 952 7274 980 12242
rect 940 7268 992 7274
rect 940 7210 992 7216
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 664 6180 716 6186
rect 664 6122 716 6128
rect 1044 5914 1072 16546
rect 1504 15706 1532 17070
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1504 13938 1532 15642
rect 1596 15502 1624 16390
rect 1688 16114 1716 16526
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1688 15026 1716 16050
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1688 14414 1716 14962
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1216 13252 1268 13258
rect 1216 13194 1268 13200
rect 1122 11656 1178 11665
rect 1122 11591 1124 11600
rect 1176 11591 1178 11600
rect 1124 11562 1176 11568
rect 1124 11348 1176 11354
rect 1124 11290 1176 11296
rect 1136 6798 1164 11290
rect 1124 6792 1176 6798
rect 1124 6734 1176 6740
rect 1032 5908 1084 5914
rect 1032 5850 1084 5856
rect 1228 5778 1256 13194
rect 1308 12980 1360 12986
rect 1308 12922 1360 12928
rect 1320 12306 1348 12922
rect 1504 12306 1532 13874
rect 1872 13002 1900 19200
rect 2042 17096 2098 17105
rect 2042 17031 2098 17040
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 14006 1992 15302
rect 1952 14000 2004 14006
rect 1952 13942 2004 13948
rect 1964 13394 1992 13942
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 13190 1992 13330
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1872 12974 1992 13002
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1308 12164 1360 12170
rect 1308 12106 1360 12112
rect 1320 7206 1348 12106
rect 1504 11762 1532 12242
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11218 1532 11698
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1504 10130 1532 11154
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1596 8090 1624 10474
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1308 7200 1360 7206
rect 1308 7142 1360 7148
rect 1216 5772 1268 5778
rect 1216 5714 1268 5720
rect 1596 5370 1624 7822
rect 1688 7478 1716 8502
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1780 6458 1808 12038
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 6662 1900 11018
rect 1964 9926 1992 12974
rect 2056 11121 2084 17031
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2042 11112 2098 11121
rect 2042 11047 2098 11056
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 7886 1992 8842
rect 2056 8090 2084 10542
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 2056 6458 2084 8026
rect 2148 7546 2176 11698
rect 2240 10810 2268 16050
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2226 10704 2282 10713
rect 2226 10639 2282 10648
rect 2240 10470 2268 10639
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2240 6662 2268 9930
rect 2332 9489 2360 14962
rect 2608 13977 2636 19200
rect 3344 19122 3372 19200
rect 3436 19122 3464 19230
rect 3344 19094 3464 19122
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16658 3004 17070
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 3528 16726 3556 16934
rect 3516 16720 3568 16726
rect 3516 16662 3568 16668
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3344 16182 3372 16458
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15570 3096 15846
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2962 15464 3018 15473
rect 2962 15399 3018 15408
rect 3056 15428 3108 15434
rect 2870 15056 2926 15065
rect 2870 14991 2926 15000
rect 2594 13968 2650 13977
rect 2594 13903 2650 13912
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2608 13462 2636 13738
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 2596 12776 2648 12782
rect 2700 12753 2728 12854
rect 2596 12718 2648 12724
rect 2686 12744 2742 12753
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2516 10713 2544 11018
rect 2502 10704 2558 10713
rect 2502 10639 2558 10648
rect 2608 10470 2636 12718
rect 2686 12679 2742 12688
rect 2700 11014 2728 12679
rect 2778 12608 2834 12617
rect 2778 12543 2834 12552
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2700 10674 2728 10950
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2424 10062 2452 10406
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9654 2452 9998
rect 2502 9888 2558 9897
rect 2502 9823 2558 9832
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2332 8634 2360 9114
rect 2424 8838 2452 9590
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2516 8786 2544 9823
rect 2700 9674 2728 10610
rect 2792 10266 2820 12543
rect 2884 12442 2912 14991
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2976 12186 3004 15399
rect 3056 15370 3108 15376
rect 3068 14278 3096 15370
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3436 14074 3464 14282
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13938 3464 14010
rect 3528 13938 3556 16662
rect 3606 16416 3662 16425
rect 3606 16351 3662 16360
rect 3620 16114 3648 16351
rect 3712 16153 3740 19230
rect 4066 19200 4122 20000
rect 4802 19200 4858 20000
rect 5538 19200 5594 20000
rect 6274 19200 6330 20000
rect 7010 19200 7066 20000
rect 7746 19200 7802 20000
rect 8482 19200 8538 20000
rect 9218 19200 9274 20000
rect 9954 19200 10010 20000
rect 10690 19200 10746 20000
rect 11426 19200 11482 20000
rect 11532 19230 11744 19258
rect 4080 17218 4108 19200
rect 3988 17190 4108 17218
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3698 16144 3754 16153
rect 3608 16108 3660 16114
rect 3698 16079 3754 16088
rect 3608 16050 3660 16056
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3620 15162 3648 15914
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15745 3740 15846
rect 3698 15736 3754 15745
rect 3698 15671 3754 15680
rect 3712 15570 3740 15671
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3804 15026 3832 16934
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3988 16538 4016 17190
rect 4344 16584 4396 16590
rect 3896 16250 3924 16526
rect 3988 16510 4108 16538
rect 4344 16526 4396 16532
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 4080 16130 4108 16510
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 3884 16108 3936 16114
rect 4080 16102 4200 16130
rect 3884 16050 3936 16056
rect 3896 15434 3924 16050
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3988 15026 4016 15846
rect 4080 15026 4108 15982
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4172 14906 4200 16102
rect 4264 15978 4292 16458
rect 4356 16425 4384 16526
rect 4436 16448 4488 16454
rect 4342 16416 4398 16425
rect 4488 16408 4660 16436
rect 4436 16390 4488 16396
rect 4342 16351 4398 16360
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4356 15858 4384 16118
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 3712 14878 4200 14906
rect 4264 15830 4384 15858
rect 3606 14240 3662 14249
rect 3606 14175 3662 14184
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 3528 13394 3556 13874
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 2884 12158 3004 12186
rect 2884 11898 2912 12158
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2870 11384 2926 11393
rect 2870 11319 2926 11328
rect 2884 11218 2912 11319
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2976 10742 3004 12038
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2976 10130 3004 10678
rect 3068 10130 3096 12718
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11558 3464 12038
rect 3528 11830 3556 12718
rect 3620 11937 3648 14175
rect 3712 12889 3740 14878
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3896 14074 3924 14554
rect 3974 14376 4030 14385
rect 3974 14311 4030 14320
rect 3988 14278 4016 14311
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 4160 14272 4212 14278
rect 4264 14260 4292 15830
rect 4448 14618 4476 15914
rect 4540 15065 4568 16186
rect 4526 15056 4582 15065
rect 4526 14991 4528 15000
rect 4580 14991 4582 15000
rect 4528 14962 4580 14968
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4344 14408 4396 14414
rect 4540 14362 4568 14962
rect 4632 14822 4660 16408
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4620 14816 4672 14822
rect 4618 14784 4620 14793
rect 4672 14784 4674 14793
rect 4618 14719 4674 14728
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4344 14350 4396 14356
rect 4212 14232 4292 14260
rect 4160 14214 4212 14220
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3804 13297 3832 13738
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3790 13288 3846 13297
rect 3790 13223 3846 13232
rect 3698 12880 3754 12889
rect 3698 12815 3754 12824
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3712 12170 3740 12650
rect 3804 12306 3832 12786
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3606 11928 3662 11937
rect 3606 11863 3662 11872
rect 3516 11824 3568 11830
rect 3896 11812 3924 13359
rect 3988 13258 4016 14214
rect 4172 14006 4200 14214
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 4172 13870 4200 13942
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4252 12912 4304 12918
rect 4356 12900 4384 14350
rect 4304 12872 4384 12900
rect 4448 14334 4568 14362
rect 4448 12900 4476 14334
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 13734 4568 14214
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4632 13190 4660 14486
rect 4724 13569 4752 16050
rect 4816 16017 4844 19200
rect 5552 17542 5580 19200
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4802 16008 4858 16017
rect 4802 15943 4858 15952
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4710 13560 4766 13569
rect 4710 13495 4766 13504
rect 4710 13424 4766 13433
rect 4710 13359 4766 13368
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4724 13025 4752 13359
rect 4710 13016 4766 13025
rect 4816 12986 4844 15846
rect 4908 15706 4936 16390
rect 5000 15978 5028 16390
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5092 15586 5120 17002
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 15978 5212 16934
rect 5448 16584 5500 16590
rect 5446 16552 5448 16561
rect 5500 16552 5502 16561
rect 5446 16487 5502 16496
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 5736 16046 5764 17138
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5172 15972 5224 15978
rect 5172 15914 5224 15920
rect 5000 15558 5120 15586
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4908 14822 4936 15098
rect 5000 15094 5028 15558
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 15162 5120 15438
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 4988 15088 5040 15094
rect 5184 15042 5212 15302
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 5540 15088 5592 15094
rect 4988 15030 5040 15036
rect 5092 15014 5212 15042
rect 5538 15056 5540 15065
rect 5592 15056 5594 15065
rect 5356 15020 5408 15026
rect 5092 14958 5120 15014
rect 5538 14991 5594 15000
rect 5356 14962 5408 14968
rect 5080 14952 5132 14958
rect 5368 14929 5396 14962
rect 5448 14952 5500 14958
rect 5080 14894 5132 14900
rect 5354 14920 5410 14929
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 13258 4936 14758
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 4710 12951 4766 12960
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4528 12912 4580 12918
rect 4448 12872 4528 12900
rect 4252 12854 4304 12860
rect 4528 12854 4580 12860
rect 4804 12776 4856 12782
rect 4710 12744 4766 12753
rect 5000 12753 5028 14418
rect 5092 13938 5120 14894
rect 5448 14894 5500 14900
rect 5354 14855 5410 14864
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 12986 5120 13738
rect 5184 13326 5212 14554
rect 5460 14550 5488 14894
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5262 14376 5318 14385
rect 5460 14346 5488 14486
rect 5552 14482 5580 14991
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5262 14311 5264 14320
rect 5316 14311 5318 14320
rect 5448 14340 5500 14346
rect 5264 14282 5316 14288
rect 5448 14282 5500 14288
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4804 12718 4856 12724
rect 4986 12744 5042 12753
rect 4710 12679 4712 12688
rect 4764 12679 4766 12688
rect 4712 12650 4764 12656
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4356 12434 4384 12582
rect 4620 12436 4672 12442
rect 4356 12406 4568 12434
rect 4342 12200 4398 12209
rect 4068 12164 4120 12170
rect 4342 12135 4398 12144
rect 4068 12106 4120 12112
rect 4080 12050 4108 12106
rect 3516 11766 3568 11772
rect 3804 11784 3924 11812
rect 3988 12022 4108 12050
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 3528 11286 3556 11766
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2962 10024 3018 10033
rect 2962 9959 3018 9968
rect 3056 9988 3108 9994
rect 2872 9716 2924 9722
rect 2596 9648 2648 9654
rect 2700 9646 2820 9674
rect 2872 9658 2924 9664
rect 2792 9602 2820 9646
rect 2596 9590 2648 9596
rect 2608 8906 2636 9590
rect 2700 9574 2820 9602
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2516 8758 2636 8786
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 7886 2360 8230
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2424 7750 2452 8570
rect 2608 8498 2636 8758
rect 2700 8566 2728 9574
rect 2780 9512 2832 9518
rect 2884 9489 2912 9658
rect 2780 9454 2832 9460
rect 2870 9480 2926 9489
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2792 8498 2820 9454
rect 2870 9415 2926 9424
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2608 8090 2636 8434
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8090 2728 8366
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 7818 2820 8434
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2332 7274 2360 7686
rect 2884 7546 2912 8842
rect 2976 8242 3004 9959
rect 3056 9930 3108 9936
rect 3068 9042 3096 9930
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9489 3464 9862
rect 3528 9586 3556 11222
rect 3620 9586 3648 11630
rect 3804 11608 3832 11784
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3712 11580 3832 11608
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3422 9480 3478 9489
rect 3478 9438 3556 9466
rect 3422 9415 3478 9424
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 3056 9036 3108 9042
rect 3528 9024 3556 9438
rect 3056 8978 3108 8984
rect 3344 8996 3556 9024
rect 3344 8634 3372 8996
rect 3514 8936 3570 8945
rect 3424 8900 3476 8906
rect 3514 8871 3570 8880
rect 3424 8842 3476 8848
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8498 3464 8842
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3436 8294 3464 8434
rect 3424 8288 3476 8294
rect 2976 8214 3096 8242
rect 3424 8230 3476 8236
rect 2962 8120 3018 8129
rect 2962 8055 3018 8064
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1582 5264 1638 5273
rect 2792 5234 2820 6831
rect 2870 6488 2926 6497
rect 2976 6474 3004 8055
rect 3068 7970 3096 8214
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 3068 7942 3188 7970
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 6798 3096 7822
rect 3160 7342 3188 7942
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2976 6446 3096 6474
rect 2870 6423 2926 6432
rect 2884 5234 2912 6423
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2976 6089 3004 6326
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 3068 5914 3096 6446
rect 3528 6322 3556 8871
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3620 5846 3648 9522
rect 3712 9217 3740 11580
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3804 9926 3832 10610
rect 3896 10033 3924 11630
rect 3988 10674 4016 12022
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3974 10568 4030 10577
rect 3974 10503 4030 10512
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3698 9208 3754 9217
rect 3698 9143 3754 9152
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3712 8430 3740 9046
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 8294 3740 8366
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3804 8022 3832 9522
rect 3896 9450 3924 9959
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3896 6866 3924 8774
rect 3988 8090 4016 10503
rect 4080 9874 4108 11494
rect 4264 10062 4292 11494
rect 4356 11370 4384 12135
rect 4540 11898 4568 12406
rect 4620 12378 4672 12384
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4448 11529 4476 11834
rect 4434 11520 4490 11529
rect 4434 11455 4490 11464
rect 4356 11342 4476 11370
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 10056 4304 10062
rect 4158 10024 4214 10033
rect 4252 9998 4304 10004
rect 4158 9959 4160 9968
rect 4212 9959 4214 9968
rect 4160 9930 4212 9936
rect 4080 9846 4200 9874
rect 4172 9654 4200 9846
rect 4160 9648 4212 9654
rect 4066 9616 4122 9625
rect 4160 9590 4212 9596
rect 4066 9551 4068 9560
rect 4120 9551 4122 9560
rect 4068 9522 4120 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4250 9480 4306 9489
rect 4172 9353 4200 9454
rect 4356 9450 4384 11222
rect 4448 10713 4476 11342
rect 4540 11150 4568 11834
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10441 4568 10610
rect 4526 10432 4582 10441
rect 4526 10367 4582 10376
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9518 4476 9862
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4250 9415 4306 9424
rect 4344 9444 4396 9450
rect 4158 9344 4214 9353
rect 4158 9279 4214 9288
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4066 8528 4122 8537
rect 4172 8498 4200 8910
rect 4264 8906 4292 9415
rect 4344 9386 4396 9392
rect 4342 9208 4398 9217
rect 4342 9143 4398 9152
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4250 8800 4306 8809
rect 4250 8735 4306 8744
rect 4066 8463 4122 8472
rect 4160 8492 4212 8498
rect 4080 8430 4108 8463
rect 4160 8434 4212 8440
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4066 7712 4122 7721
rect 4066 7647 4122 7656
rect 4080 7342 4108 7647
rect 4068 7336 4120 7342
rect 3974 7304 4030 7313
rect 4068 7278 4120 7284
rect 3974 7239 4030 7248
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3988 6730 4016 7239
rect 4172 6934 4200 8434
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4264 6866 4292 8735
rect 4356 8498 4384 9143
rect 4540 9110 4568 10202
rect 4632 9926 4660 12378
rect 4816 12102 4844 12718
rect 4986 12679 5042 12688
rect 5276 12345 5304 13942
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5368 13190 5396 13874
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5644 13394 5672 13806
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 5388 13019 5696 13028
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5262 12336 5318 12345
rect 5262 12271 5318 12280
rect 4986 12200 5042 12209
rect 4986 12135 4988 12144
rect 5040 12135 5042 12144
rect 5080 12164 5132 12170
rect 4988 12106 5040 12112
rect 5080 12106 5132 12112
rect 4804 12096 4856 12102
rect 5092 12050 5120 12106
rect 5644 12084 5672 12650
rect 5736 12434 5764 15982
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5828 14890 5856 15302
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5920 14550 5948 16934
rect 6012 16697 6040 16934
rect 5998 16688 6054 16697
rect 5998 16623 6054 16632
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6012 15337 6040 16186
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 5998 15328 6054 15337
rect 5998 15263 6054 15272
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 6012 14414 6040 15030
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 13530 5856 14214
rect 5906 13832 5962 13841
rect 5906 13767 5962 13776
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5828 13025 5856 13466
rect 5920 13274 5948 13767
rect 6012 13530 6040 14350
rect 6104 14278 6132 15914
rect 6196 14521 6224 16458
rect 6182 14512 6238 14521
rect 6182 14447 6238 14456
rect 6288 14464 6316 19200
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17270 6592 17546
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6564 16522 6592 17206
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16182 6592 16458
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6288 14436 6408 14464
rect 6274 14376 6330 14385
rect 6274 14311 6330 14320
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5920 13246 6132 13274
rect 6000 13184 6052 13190
rect 5920 13144 6000 13172
rect 5814 13016 5870 13025
rect 5814 12951 5870 12960
rect 5736 12406 5856 12434
rect 5644 12056 5764 12084
rect 4804 12038 4856 12044
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4724 10062 4752 11698
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4632 9450 4660 9590
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4632 8906 4660 9386
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3988 5914 4016 6666
rect 4356 6458 4384 8434
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3976 5704 4028 5710
rect 3974 5672 3976 5681
rect 4028 5672 4030 5681
rect 4448 5642 4476 8298
rect 4632 8294 4660 8842
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4724 8090 4752 9998
rect 4816 8974 4844 12038
rect 5000 12022 5120 12050
rect 5000 11830 5028 12022
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 5736 11830 5764 12056
rect 4988 11824 5040 11830
rect 5724 11824 5776 11830
rect 4988 11766 5040 11772
rect 5078 11792 5134 11801
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4908 9654 4936 11698
rect 5000 10062 5028 11766
rect 5724 11766 5776 11772
rect 5078 11727 5134 11736
rect 5264 11756 5316 11762
rect 5092 11694 5120 11727
rect 5264 11698 5316 11704
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5276 11506 5304 11698
rect 5354 11656 5410 11665
rect 5354 11591 5356 11600
rect 5408 11591 5410 11600
rect 5356 11562 5408 11568
rect 5724 11552 5776 11558
rect 5092 11150 5120 11494
rect 5276 11478 5396 11506
rect 5724 11494 5776 11500
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5184 11150 5212 11222
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5080 11008 5132 11014
rect 5172 11008 5224 11014
rect 5080 10950 5132 10956
rect 5170 10976 5172 10985
rect 5224 10976 5226 10985
rect 5092 10266 5120 10950
rect 5170 10911 5226 10920
rect 5170 10432 5226 10441
rect 5170 10367 5226 10376
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5000 9178 5028 9454
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 5092 7546 5120 10066
rect 5184 8294 5212 10367
rect 5276 10266 5304 11290
rect 5368 11286 5396 11478
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 5538 10704 5594 10713
rect 5538 10639 5540 10648
rect 5592 10639 5594 10648
rect 5540 10610 5592 10616
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 10146 5396 10542
rect 5552 10266 5580 10610
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5276 10118 5396 10146
rect 5276 9926 5304 10118
rect 5446 10024 5502 10033
rect 5446 9959 5448 9968
rect 5500 9959 5502 9968
rect 5448 9930 5500 9936
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9353 5304 9862
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 5736 9654 5764 11494
rect 5724 9648 5776 9654
rect 5630 9616 5686 9625
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5448 9580 5500 9586
rect 5724 9590 5776 9596
rect 5630 9551 5686 9560
rect 5448 9522 5500 9528
rect 5262 9344 5318 9353
rect 5262 9279 5318 9288
rect 5368 8974 5396 9522
rect 5460 9042 5488 9522
rect 5538 9208 5594 9217
rect 5538 9143 5540 9152
rect 5592 9143 5594 9152
rect 5540 9114 5592 9120
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5644 8820 5672 9551
rect 5644 8792 5764 8820
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 5736 8498 5764 8792
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5262 8120 5318 8129
rect 5262 8055 5264 8064
rect 5316 8055 5318 8064
rect 5264 8026 5316 8032
rect 5644 7954 5672 8230
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 3974 5607 4030 5616
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4540 5302 4568 6802
rect 5736 6798 5764 8434
rect 5828 7546 5856 12406
rect 5920 11218 5948 13144
rect 6000 13126 6052 13132
rect 5998 13016 6054 13025
rect 5998 12951 6054 12960
rect 6012 12238 6040 12951
rect 6104 12782 6132 13246
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5920 10538 5948 11018
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5920 8906 5948 9658
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5814 7440 5870 7449
rect 5814 7375 5816 7384
rect 5868 7375 5870 7384
rect 5816 7346 5868 7352
rect 5828 7002 5856 7346
rect 5920 7274 5948 7822
rect 6012 7478 6040 12174
rect 6104 11370 6132 12718
rect 6196 12170 6224 13194
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6288 11558 6316 14311
rect 6380 12458 6408 14436
rect 6472 14090 6500 15506
rect 6656 15366 6684 16594
rect 6840 16590 6868 16934
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6748 15178 6776 15438
rect 6656 15150 6776 15178
rect 6472 14062 6592 14090
rect 6460 13864 6512 13870
rect 6458 13832 6460 13841
rect 6512 13832 6514 13841
rect 6458 13767 6514 13776
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6472 12714 6500 12854
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6380 12430 6500 12458
rect 6564 12442 6592 14062
rect 6656 13938 6684 15150
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6472 12220 6500 12430
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6656 12374 6684 13466
rect 6748 12374 6776 14758
rect 6840 13530 6868 15914
rect 6932 15434 6960 16186
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 14414 6960 15370
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6932 13410 6960 13942
rect 6840 13382 6960 13410
rect 6840 12442 6868 13382
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6828 12232 6880 12238
rect 6472 12192 6684 12220
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6104 11342 6316 11370
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 1582 5199 1638 5208
rect 2780 5228 2832 5234
rect 1596 4146 1624 5199
rect 2780 5170 2832 5176
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 6104 4622 6132 9862
rect 6196 9674 6224 11154
rect 6288 11150 6316 11342
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6196 9646 6316 9674
rect 6182 9072 6238 9081
rect 6182 9007 6238 9016
rect 6196 8974 6224 9007
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6196 7546 6224 8910
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7206 6316 9646
rect 6380 7342 6408 12106
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6472 6730 6500 11698
rect 6564 10674 6592 11834
rect 6656 11150 6684 12192
rect 6828 12174 6880 12180
rect 6840 11354 6868 12174
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6748 10266 6776 11018
rect 6932 10810 6960 12582
rect 7024 11762 7052 19200
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 15994 7144 17478
rect 7760 17082 7788 19200
rect 7760 17054 7972 17082
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 16289 7236 16934
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 7288 16584 7340 16590
rect 7340 16532 7512 16538
rect 7288 16526 7512 16532
rect 7300 16510 7512 16526
rect 7288 16448 7340 16454
rect 7340 16408 7420 16436
rect 7288 16390 7340 16396
rect 7194 16280 7250 16289
rect 7194 16215 7250 16224
rect 7208 16114 7236 16215
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7116 15966 7236 15994
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15706 7144 15846
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7208 15552 7236 15966
rect 7300 15638 7328 16118
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7116 15524 7236 15552
rect 7116 13784 7144 15524
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 14346 7236 15302
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14618 7328 15030
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7116 13756 7328 13784
rect 7194 13696 7250 13705
rect 7194 13631 7250 13640
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7010 11520 7066 11529
rect 7010 11455 7066 11464
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6564 8022 6592 10202
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9489 6684 9998
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6826 9208 6882 9217
rect 7024 9178 7052 11455
rect 6826 9143 6828 9152
rect 6880 9143 6882 9152
rect 7012 9172 7064 9178
rect 6828 9114 6880 9120
rect 7012 9114 7064 9120
rect 7116 8974 7144 13262
rect 7208 11200 7236 13631
rect 7300 12356 7328 13756
rect 7392 13258 7420 16408
rect 7484 15065 7512 16510
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7668 16182 7696 16390
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7838 16008 7894 16017
rect 7838 15943 7894 15952
rect 7852 15910 7880 15943
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7470 15056 7526 15065
rect 7470 14991 7526 15000
rect 7576 14890 7604 15642
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7748 15496 7800 15502
rect 7746 15464 7748 15473
rect 7800 15464 7802 15473
rect 7746 15399 7802 15408
rect 7852 15201 7880 15574
rect 7838 15192 7894 15201
rect 7838 15127 7894 15136
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 13530 7512 14758
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7576 14362 7604 14486
rect 7576 14346 7880 14362
rect 7576 14340 7892 14346
rect 7576 14334 7840 14340
rect 7840 14282 7892 14288
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7852 13870 7880 14010
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7668 13433 7696 13466
rect 7748 13456 7800 13462
rect 7654 13424 7710 13433
rect 7748 13398 7800 13404
rect 7654 13359 7710 13368
rect 7760 13326 7788 13398
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12646 7512 13126
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7576 12714 7604 12922
rect 7656 12776 7708 12782
rect 7654 12744 7656 12753
rect 7708 12744 7710 12753
rect 7564 12708 7616 12714
rect 7654 12679 7710 12688
rect 7564 12650 7616 12656
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 7300 12328 7420 12356
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7300 11354 7328 11630
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7208 11172 7328 11200
rect 7194 11112 7250 11121
rect 7194 11047 7250 11056
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7208 8820 7236 11047
rect 7300 10606 7328 11172
rect 7392 10674 7420 12328
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7484 11354 7512 12106
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11830 7696 12038
rect 7760 11898 7788 12174
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7944 11762 7972 17054
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8206 16280 8262 16289
rect 8206 16215 8262 16224
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8036 15638 8064 16118
rect 8114 15872 8170 15881
rect 8114 15807 8170 15816
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8036 14958 8064 15574
rect 8128 15434 8156 15807
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8114 15192 8170 15201
rect 8114 15127 8170 15136
rect 8128 15094 8156 15127
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8128 14958 8156 15030
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8022 14512 8078 14521
rect 8220 14482 8248 16215
rect 8312 16182 8340 16390
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15881 8340 15982
rect 8298 15872 8354 15881
rect 8298 15807 8354 15816
rect 8404 15638 8432 16390
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8312 14929 8340 15030
rect 8298 14920 8354 14929
rect 8298 14855 8354 14864
rect 8404 14618 8432 15574
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8022 14447 8078 14456
rect 8208 14476 8260 14482
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9722 7604 9998
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7116 8792 7236 8820
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 7116 7886 7144 8792
rect 7944 8634 7972 11562
rect 8036 10266 8064 14447
rect 8208 14418 8260 14424
rect 8220 13938 8248 14418
rect 8496 14090 8524 19200
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17134 8616 17614
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8680 16114 8708 16458
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8666 16008 8722 16017
rect 8666 15943 8722 15952
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8404 14062 8524 14090
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 11286 8156 13806
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13394 8248 13670
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8206 13288 8262 13297
rect 8206 13223 8262 13232
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10606 8156 11086
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9110 8064 9998
rect 8220 9586 8248 13223
rect 8404 12434 8432 14062
rect 8588 14006 8616 14758
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8496 13870 8524 13942
rect 8484 13864 8536 13870
rect 8482 13832 8484 13841
rect 8536 13832 8538 13841
rect 8482 13767 8538 13776
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13258 8524 13670
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8312 12406 8432 12434
rect 8312 12238 8340 12406
rect 8496 12306 8524 13194
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8588 12238 8616 13262
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8680 11762 8708 15943
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 15434 8800 15574
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 12986 8800 15098
rect 8864 14822 8892 16050
rect 8956 15570 8984 16526
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14414 8892 14758
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 14006 8892 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8864 12850 8892 13942
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8956 12238 8984 15302
rect 9048 12442 9076 16050
rect 9140 15706 9168 17138
rect 9232 15706 9260 19200
rect 9968 17746 9996 19200
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17338 9720 17478
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9324 15473 9352 17138
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16114 9628 16390
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9310 15464 9366 15473
rect 9310 15399 9366 15408
rect 9324 15366 9352 15399
rect 9312 15360 9364 15366
rect 9218 15328 9274 15337
rect 9312 15302 9364 15308
rect 9218 15263 9274 15272
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 14074 9168 14350
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 12850 9168 13874
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9128 12368 9180 12374
rect 9126 12336 9128 12345
rect 9180 12336 9182 12345
rect 9126 12271 9182 12280
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8666 10704 8722 10713
rect 9232 10674 9260 15263
rect 9324 13326 9352 15302
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9416 14278 9444 15098
rect 9508 14414 9536 15846
rect 9600 14958 9628 16050
rect 9692 15502 9720 17138
rect 10520 17134 10548 17614
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 17338 10640 17546
rect 10704 17542 10732 19200
rect 11440 19122 11468 19200
rect 11532 19122 11560 19230
rect 11440 19094 11560 19122
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9600 14346 9628 14894
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9692 14074 9720 14962
rect 9876 14482 9904 15030
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9508 13462 9536 13738
rect 9496 13456 9548 13462
rect 9402 13424 9458 13433
rect 9496 13398 9548 13404
rect 9402 13359 9404 13368
rect 9456 13359 9458 13368
rect 9404 13330 9456 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9588 13184 9640 13190
rect 9784 13172 9812 13738
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 13297 9904 13330
rect 9862 13288 9918 13297
rect 9862 13223 9918 13232
rect 9968 13190 9996 14010
rect 10152 13734 10180 14010
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10244 13512 10272 16458
rect 10336 14618 10364 17070
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10060 13484 10272 13512
rect 9588 13126 9640 13132
rect 9692 13144 9812 13172
rect 9956 13184 10008 13190
rect 9310 12880 9366 12889
rect 9600 12850 9628 13126
rect 9692 12968 9720 13144
rect 10060 13172 10088 13484
rect 10060 13144 10272 13172
rect 9956 13126 10008 13132
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 10244 12986 10272 13144
rect 10232 12980 10284 12986
rect 9692 12940 9812 12968
rect 9678 12880 9734 12889
rect 9310 12815 9366 12824
rect 9496 12844 9548 12850
rect 9324 11150 9352 12815
rect 9496 12786 9548 12792
rect 9588 12844 9640 12850
rect 9678 12815 9734 12824
rect 9588 12786 9640 12792
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9416 12646 9444 12718
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9508 12434 9536 12786
rect 9508 12406 9628 12434
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9416 11626 9444 11834
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9600 11778 9628 12406
rect 9692 11898 9720 12815
rect 9784 12442 9812 12940
rect 10232 12922 10284 12928
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12481 10180 12582
rect 10138 12472 10194 12481
rect 9772 12436 9824 12442
rect 10138 12407 10194 12416
rect 9772 12378 9824 12384
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 10060 12238 10088 12271
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10230 12200 10286 12209
rect 10230 12135 10286 12144
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 10244 11898 10272 12135
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9508 11218 9536 11766
rect 9600 11750 9720 11778
rect 9692 11354 9720 11750
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8666 10639 8668 10648
rect 8720 10639 8722 10648
rect 9220 10668 9272 10674
rect 8668 10610 8720 10616
rect 9220 10610 9272 10616
rect 9126 10296 9182 10305
rect 9324 10266 9352 11086
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 10336 10810 10364 14418
rect 10428 13802 10456 17002
rect 10520 16590 10548 17070
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10520 15201 10548 15574
rect 10506 15192 10562 15201
rect 10506 15127 10562 15136
rect 10506 14920 10562 14929
rect 10506 14855 10508 14864
rect 10560 14855 10562 14864
rect 10508 14826 10560 14832
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 14260 10548 14554
rect 10612 14414 10640 15846
rect 10704 15502 10732 16526
rect 10796 16114 10824 17206
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16250 11008 16390
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15496 10744 15502
rect 10690 15464 10692 15473
rect 10744 15464 10746 15473
rect 10690 15399 10746 15408
rect 10692 15360 10744 15366
rect 10690 15328 10692 15337
rect 10744 15328 10746 15337
rect 10690 15263 10746 15272
rect 10796 15162 10824 16050
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10782 15056 10838 15065
rect 10782 14991 10838 15000
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10520 14232 10640 14260
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10414 13424 10470 13433
rect 10414 13359 10470 13368
rect 10428 13326 10456 13359
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10506 12472 10562 12481
rect 10506 12407 10562 12416
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10428 11898 10456 12242
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9126 10231 9128 10240
rect 9180 10231 9182 10240
rect 9312 10260 9364 10266
rect 9128 10202 9180 10208
rect 9312 10202 9364 10208
rect 8666 9616 8722 9625
rect 8208 9580 8260 9586
rect 8666 9551 8668 9560
rect 8208 9522 8260 9528
rect 8720 9551 8722 9560
rect 9126 9616 9182 9625
rect 9126 9551 9128 9560
rect 8668 9522 8720 9528
rect 9180 9551 9182 9560
rect 9128 9522 9180 9528
rect 8114 9480 8170 9489
rect 8114 9415 8170 9424
rect 8128 9178 8156 9415
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7194 8528 7250 8537
rect 7194 8463 7196 8472
rect 7248 8463 7250 8472
rect 7196 8434 7248 8440
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7116 7546 7144 7822
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 8496 6866 8524 9318
rect 8680 9178 8708 9522
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 9600 8090 9628 10610
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9654 9720 9998
rect 10520 9994 10548 12407
rect 10612 11830 10640 14232
rect 10704 12102 10732 14826
rect 10796 12850 10824 14991
rect 10888 12986 10916 15370
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10980 15094 11008 15302
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10980 12850 11008 13398
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11072 12442 11100 17138
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11164 16250 11192 16730
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 15570 11284 17274
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11164 12850 11192 14758
rect 11256 14618 11284 14962
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11256 13938 11284 14214
rect 11348 14074 11376 14214
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11256 13326 11284 13874
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10888 11898 10916 12310
rect 11256 12238 11284 12718
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10600 11824 10652 11830
rect 11164 11801 11192 12174
rect 10600 11766 10652 11772
rect 11150 11792 11206 11801
rect 10876 11756 10928 11762
rect 11150 11727 11206 11736
rect 10876 11698 10928 11704
rect 10888 11558 10916 11698
rect 11440 11626 11468 16458
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 14006 11560 16050
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 13326 11560 13466
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11624 12986 11652 16730
rect 11716 16590 11744 19230
rect 12162 19200 12218 20000
rect 12898 19200 12954 20000
rect 13634 19200 13690 20000
rect 14370 19200 14426 20000
rect 15106 19200 15162 20000
rect 15842 19200 15898 20000
rect 16578 19200 16634 20000
rect 16684 19230 16896 19258
rect 12176 16980 12204 19200
rect 11992 16952 12204 16980
rect 11992 16946 12020 16952
rect 11972 16918 12020 16946
rect 11972 16810 12000 16918
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 11972 16782 12020 16810
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 15978 11836 16390
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 14958 11744 15846
rect 11808 15434 11836 15914
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11716 14074 11744 14282
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11808 13870 11836 14758
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11900 13530 11928 15982
rect 11992 15858 12020 16782
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12360 16522 12388 16730
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 16046 12296 16118
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 11972 15830 12020 15858
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 11972 15722 12000 15830
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 11972 15694 12020 15722
rect 11992 15026 12020 15694
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 15094 12112 15506
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12176 14929 12204 15574
rect 12452 15434 12480 15846
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12438 15192 12494 15201
rect 12438 15127 12494 15136
rect 12162 14920 12218 14929
rect 12162 14855 12218 14864
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 12452 14618 12480 15127
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14278 12572 15302
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12636 13734 12664 16730
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12728 15570 12756 15642
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 12728 13546 12756 15302
rect 12820 15162 12848 16390
rect 12912 16130 12940 19200
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 12912 16102 13032 16130
rect 13096 16114 13124 16662
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12912 14346 12940 15982
rect 13004 15570 13032 16102
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13082 16008 13138 16017
rect 13082 15943 13138 15952
rect 13176 15972 13228 15978
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13004 15337 13032 15370
rect 12990 15328 13046 15337
rect 12990 15263 13046 15272
rect 13096 14550 13124 15943
rect 13176 15914 13228 15920
rect 13188 15094 13216 15914
rect 13280 15706 13308 16458
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13280 15502 13308 15642
rect 13358 15600 13414 15609
rect 13358 15535 13414 15544
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14550 13216 14758
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12898 13832 12954 13841
rect 12898 13767 12954 13776
rect 11888 13524 11940 13530
rect 12728 13518 12848 13546
rect 11888 13466 11940 13472
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11808 12442 11836 12650
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 12820 12306 12848 13518
rect 12912 13326 12940 13767
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 13096 12434 13124 14350
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13004 12406 13124 12434
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 13004 12170 13032 12406
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 11702 11792 11758 11801
rect 11702 11727 11704 11736
rect 11756 11727 11758 11736
rect 11704 11698 11756 11704
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 11060 11280 11112 11286
rect 11058 11248 11060 11257
rect 11112 11248 11114 11257
rect 11058 11183 11114 11192
rect 13280 11014 13308 13330
rect 13372 13190 13400 15535
rect 13464 14482 13492 16118
rect 13556 15638 13584 17682
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13648 15450 13676 19200
rect 14384 17626 14412 19200
rect 14200 17598 14412 17626
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 17202 13768 17478
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13648 15422 13860 15450
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13542 15056 13598 15065
rect 13542 14991 13598 15000
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13464 12986 13492 14418
rect 13556 13394 13584 14991
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13648 11354 13676 15302
rect 13740 13938 13768 15302
rect 13832 14618 13860 15422
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13818 14376 13874 14385
rect 13818 14311 13874 14320
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13832 12850 13860 14311
rect 13924 14074 13952 16458
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13910 13560 13966 13569
rect 13910 13495 13966 13504
rect 13924 12918 13952 13495
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 14016 12646 14044 15574
rect 14108 15434 14136 15982
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14108 11898 14136 15370
rect 14200 13938 14228 17598
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16590 14320 16934
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14384 15609 14412 16118
rect 14370 15600 14426 15609
rect 14568 15570 14596 16186
rect 14370 15535 14426 15544
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14346 15088 14398 15094
rect 14398 15036 14412 15076
rect 14346 15030 14412 15036
rect 14384 14346 14412 15030
rect 14568 14890 14596 15098
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14660 14822 14688 16390
rect 14936 16046 14964 17070
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14924 16040 14976 16046
rect 14922 16008 14924 16017
rect 14976 16008 14978 16017
rect 14922 15943 14978 15952
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14292 13818 14320 14010
rect 14370 13968 14426 13977
rect 14370 13903 14426 13912
rect 14384 13870 14412 13903
rect 14200 13790 14320 13818
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13726 11792 13782 11801
rect 13726 11727 13728 11736
rect 13780 11727 13782 11736
rect 13728 11698 13780 11704
rect 14200 11354 14228 13790
rect 14556 13728 14608 13734
rect 14554 13696 14556 13705
rect 14608 13696 14610 13705
rect 14554 13631 14610 13640
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 14660 12850 14688 14010
rect 14752 13394 14780 15846
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14462 11384 14518 11393
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14188 11348 14240 11354
rect 14462 11319 14518 11328
rect 14188 11290 14240 11296
rect 14476 11286 14504 11319
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 14660 9450 14688 11698
rect 14752 11694 14780 12854
rect 14844 12730 14872 15642
rect 14936 12850 14964 15846
rect 15028 15706 15056 16526
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15016 15496 15068 15502
rect 15014 15464 15016 15473
rect 15068 15464 15070 15473
rect 15014 15399 15070 15408
rect 15120 14906 15148 19200
rect 15856 17218 15884 19200
rect 16592 19122 16620 19200
rect 16684 19122 16712 19230
rect 16592 19094 16712 19122
rect 16026 19000 16082 19009
rect 16026 18935 16082 18944
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15764 17190 15884 17218
rect 15028 14878 15148 14906
rect 15028 14770 15056 14878
rect 15028 14742 15148 14770
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14844 12702 14964 12730
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 11762 14872 12582
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14936 11286 14964 12702
rect 15028 12442 15056 14554
rect 15120 13326 15148 14742
rect 15212 14618 15240 17138
rect 15290 16552 15346 16561
rect 15290 16487 15292 16496
rect 15344 16487 15346 16496
rect 15292 16458 15344 16464
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15396 15706 15424 16118
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15292 15632 15344 15638
rect 15292 15574 15344 15580
rect 15658 15600 15714 15609
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 14113 15240 14282
rect 15198 14104 15254 14113
rect 15198 14039 15254 14048
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15028 11830 15056 12106
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 15120 10810 15148 13262
rect 15212 13190 15240 13942
rect 15304 13705 15332 15574
rect 15658 15535 15714 15544
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 14618 15424 14758
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15396 14414 15424 14554
rect 15580 14414 15608 14894
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15290 13696 15346 13705
rect 15290 13631 15346 13640
rect 15304 13326 15332 13631
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15200 13184 15252 13190
rect 15396 13138 15424 14350
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15488 13705 15516 13738
rect 15474 13696 15530 13705
rect 15474 13631 15530 13640
rect 15200 13126 15252 13132
rect 15304 13110 15424 13138
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15212 9518 15240 12718
rect 15304 12238 15332 13110
rect 15382 13016 15438 13025
rect 15382 12951 15438 12960
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 11762 15332 12174
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15396 10266 15424 12951
rect 15474 12880 15530 12889
rect 15474 12815 15530 12824
rect 15488 12714 15516 12815
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15488 11898 15516 12543
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15580 10198 15608 14350
rect 15672 13433 15700 15535
rect 15764 15366 15792 17190
rect 15842 17096 15898 17105
rect 15842 17031 15898 17040
rect 15856 16794 15884 17031
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15948 15706 15976 15982
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15948 15162 15976 15438
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15658 13424 15714 13433
rect 15658 13359 15714 13368
rect 15764 13326 15792 14962
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15856 14482 15884 14758
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15842 14240 15898 14249
rect 15842 14175 15898 14184
rect 15752 13320 15804 13326
rect 15658 13288 15714 13297
rect 15752 13262 15804 13268
rect 15658 13223 15714 13232
rect 15672 12850 15700 13223
rect 15750 13152 15806 13161
rect 15750 13087 15806 13096
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15764 10674 15792 13087
rect 15856 12306 15884 14175
rect 15948 13938 15976 15098
rect 16040 15065 16068 18935
rect 16394 17776 16450 17785
rect 16394 17711 16450 17720
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16026 15056 16082 15065
rect 16026 14991 16082 15000
rect 16026 14920 16082 14929
rect 16026 14855 16082 14864
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16040 13682 16068 14855
rect 15948 13654 16068 13682
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15948 11762 15976 13654
rect 16026 13424 16082 13433
rect 16026 13359 16082 13368
rect 16040 12306 16068 13359
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 16132 11354 16160 16458
rect 16224 16017 16252 16526
rect 16316 16114 16344 16934
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16210 16008 16266 16017
rect 16210 15943 16266 15952
rect 16224 15502 16252 15943
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16316 15094 16344 16050
rect 16304 15088 16356 15094
rect 16408 15065 16436 17711
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 16868 15910 16896 19230
rect 17314 19200 17370 20000
rect 17420 19230 17632 19258
rect 17328 19122 17356 19200
rect 17420 19122 17448 19230
rect 17328 19094 17448 19122
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16960 16114 16988 17070
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17144 16590 17172 16934
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 16960 15502 16988 16050
rect 16948 15496 17000 15502
rect 17144 15473 17172 16526
rect 17130 15464 17186 15473
rect 16948 15438 17000 15444
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16304 15030 16356 15036
rect 16394 15056 16450 15065
rect 16212 15020 16264 15026
rect 16394 14991 16450 15000
rect 16212 14962 16264 14968
rect 16224 14793 16252 14962
rect 16396 14816 16448 14822
rect 16210 14784 16266 14793
rect 16396 14758 16448 14764
rect 16210 14719 16266 14728
rect 16224 14396 16252 14719
rect 16304 14408 16356 14414
rect 16224 14368 16304 14396
rect 16304 14350 16356 14356
rect 16212 14272 16264 14278
rect 16210 14240 16212 14249
rect 16264 14240 16266 14249
rect 16210 14175 16266 14184
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16224 13705 16252 13942
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16210 13696 16266 13705
rect 16210 13631 16266 13640
rect 16224 13190 16252 13631
rect 16316 13326 16344 13806
rect 16408 13326 16436 14758
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 16868 14498 16896 15370
rect 16960 14958 16988 15438
rect 17052 15422 17130 15450
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14618 16988 14894
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16776 14470 16896 14498
rect 16486 14376 16542 14385
rect 16486 14311 16542 14320
rect 16500 14006 16528 14311
rect 16776 14278 16804 14470
rect 17052 14385 17080 15422
rect 17130 15399 17186 15408
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17038 14376 17094 14385
rect 17038 14311 17094 14320
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16486 13832 16542 13841
rect 16592 13818 16620 14010
rect 16542 13790 16620 13818
rect 16670 13832 16726 13841
rect 16486 13767 16542 13776
rect 16776 13802 16804 14214
rect 16946 14104 17002 14113
rect 16946 14039 17002 14048
rect 16960 14006 16988 14039
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16946 13832 17002 13841
rect 16670 13767 16726 13776
rect 16764 13796 16816 13802
rect 16684 13734 16712 13767
rect 16764 13738 16816 13744
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16868 13138 16896 13806
rect 16946 13767 17002 13776
rect 16960 13530 16988 13767
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17052 13326 17080 14214
rect 17144 13394 17172 14486
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 16868 13110 17080 13138
rect 16946 12880 17002 12889
rect 16396 12844 16448 12850
rect 16946 12815 17002 12824
rect 16396 12786 16448 12792
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16302 12744 16358 12753
rect 16224 12594 16252 12718
rect 16302 12679 16304 12688
rect 16356 12679 16358 12688
rect 16304 12650 16356 12656
rect 16224 12566 16344 12594
rect 16210 12472 16266 12481
rect 16210 12407 16266 12416
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 16224 10266 16252 12407
rect 16316 12238 16344 12566
rect 16408 12374 16436 12786
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11150 16436 12038
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16868 10674 16896 12582
rect 16960 12442 16988 12815
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17052 12170 17080 13110
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17144 11354 17172 13194
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 17144 9178 17172 11154
rect 17236 10810 17264 15370
rect 17328 13530 17356 16594
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17420 16182 17448 16526
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17420 14006 17448 15098
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17420 12918 17448 13806
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17420 12306 17448 12854
rect 17512 12442 17540 14554
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17328 11354 17356 12106
rect 17420 11898 17448 12106
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17498 11656 17554 11665
rect 17498 11591 17500 11600
rect 17552 11591 17554 11600
rect 17500 11562 17552 11568
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17420 10266 17448 11018
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17604 10062 17632 19230
rect 18050 19200 18106 20000
rect 18786 19200 18842 20000
rect 19168 19230 19472 19258
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 15502 17816 16526
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17682 14512 17738 14521
rect 17682 14447 17738 14456
rect 17696 11286 17724 14447
rect 17788 12850 17816 15030
rect 17880 12986 17908 15642
rect 17972 13569 18000 17138
rect 18064 15910 18092 19200
rect 18800 17542 18828 19200
rect 19062 18184 19118 18193
rect 19062 18119 19118 18128
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18340 16250 18368 16526
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18602 16144 18658 16153
rect 18602 16079 18658 16088
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 18064 15026 18092 15574
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18064 14362 18092 14962
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18156 14482 18184 14758
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18236 14408 18288 14414
rect 18064 14346 18184 14362
rect 18236 14350 18288 14356
rect 18064 14340 18196 14346
rect 18064 14334 18144 14340
rect 18144 14282 18196 14288
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17958 13560 18014 13569
rect 17958 13495 18014 13504
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17972 11898 18000 12650
rect 18064 12442 18092 14214
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18156 13462 18184 14010
rect 18248 13734 18276 14350
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18234 13560 18290 13569
rect 18234 13495 18290 13504
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 18156 12986 18184 13398
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17958 11792 18014 11801
rect 17958 11727 17960 11736
rect 18012 11727 18014 11736
rect 17960 11698 18012 11704
rect 18052 11688 18104 11694
rect 18156 11676 18184 12922
rect 18104 11648 18184 11676
rect 18052 11630 18104 11636
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17696 10713 17724 11086
rect 17682 10704 17738 10713
rect 17682 10639 17738 10648
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 17604 8634 17632 9998
rect 17696 9722 17724 10639
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17880 9110 17908 11086
rect 18248 10538 18276 13495
rect 18340 12986 18368 14214
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18340 11830 18368 12650
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18326 11248 18382 11257
rect 18326 11183 18382 11192
rect 18340 10674 18368 11183
rect 18432 10742 18460 15370
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18524 13190 18552 13738
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12714 18552 13126
rect 18616 12730 18644 16079
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 13530 18736 13670
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 18512 12708 18564 12714
rect 18616 12702 18828 12730
rect 18512 12650 18564 12656
rect 18800 12458 18828 12702
rect 18616 12430 18828 12458
rect 18510 11792 18566 11801
rect 18510 11727 18566 11736
rect 18524 11150 18552 11727
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18616 10606 18644 12430
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18326 10432 18382 10441
rect 18326 10367 18382 10376
rect 18340 10266 18368 10367
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18326 10024 18382 10033
rect 18326 9959 18382 9968
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17972 9042 18000 9590
rect 18340 9586 18368 9959
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 19076 9654 19104 18119
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 19168 9518 19196 19230
rect 19444 19122 19472 19230
rect 19522 19200 19578 20000
rect 19536 19122 19564 19200
rect 19444 19094 19564 19122
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 12374 19288 15846
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19444 11898 19472 17478
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 18326 9208 18382 9217
rect 18326 9143 18328 9152
rect 18380 9143 18382 9152
rect 18328 9114 18380 9120
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 19154 8800 19210 8809
rect 18705 8732 19013 8741
rect 19154 8735 19210 8744
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 19168 8498 19196 8735
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 18326 7984 18382 7993
rect 18326 7919 18328 7928
rect 18380 7919 18382 7928
rect 18328 7890 18380 7896
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 18326 7440 18382 7449
rect 18326 7375 18328 7384
rect 18380 7375 18382 7384
rect 18328 7346 18380 7352
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 18328 6792 18380 6798
rect 18326 6760 18328 6769
rect 18380 6760 18382 6769
rect 6460 6724 6512 6730
rect 18326 6695 18382 6704
rect 6460 6666 6512 6672
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 18326 6352 18382 6361
rect 18326 6287 18328 6296
rect 18380 6287 18382 6296
rect 18328 6258 18380 6264
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 18328 5704 18380 5710
rect 18326 5672 18328 5681
rect 18380 5672 18382 5681
rect 18326 5607 18382 5616
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 18326 5128 18382 5137
rect 18326 5063 18328 5072
rect 18380 5063 18382 5072
rect 18328 5034 18380 5040
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 1676 4480 1728 4486
rect 1674 4448 1676 4457
rect 1728 4448 1730 4457
rect 1674 4383 1730 4392
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 19168 4321 19196 4558
rect 19154 4312 19210 4321
rect 19154 4247 19210 4256
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1596 3738 1624 3975
rect 18328 3936 18380 3942
rect 18326 3904 18328 3913
rect 18380 3904 18382 3913
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 16486 3836 16794 3845
rect 18326 3839 18382 3848
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 1582 3224 1638 3233
rect 5388 3227 5696 3236
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 1582 3159 1638 3168
rect 1596 3058 1624 3159
rect 18340 3097 18368 3470
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 18326 3088 18382 3097
rect 1584 3052 1636 3058
rect 18326 3023 18382 3032
rect 1584 2994 1636 3000
rect 18328 2848 18380 2854
rect 1582 2816 1638 2825
rect 18328 2790 18380 2796
rect 1582 2751 1638 2760
rect 1596 2650 1624 2751
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 18340 2689 18368 2790
rect 18326 2680 18382 2689
rect 1584 2644 1636 2650
rect 18326 2615 18382 2624
rect 1584 2586 1636 2592
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 2240 2009 2268 2382
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 2884 1601 2912 2382
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 17696 1465 17724 2382
rect 18340 1873 18368 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 17682 1456 17738 1465
rect 17682 1391 17738 1400
<< via2 >>
rect 386 18536 442 18592
rect 1122 11620 1178 11656
rect 1122 11600 1124 11620
rect 1124 11600 1176 11620
rect 1176 11600 1178 11620
rect 2042 17040 2098 17096
rect 2042 11056 2098 11112
rect 2226 10648 2282 10704
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 2962 15408 3018 15464
rect 2870 15000 2926 15056
rect 2594 13912 2650 13968
rect 2502 10648 2558 10704
rect 2686 12688 2742 12744
rect 2778 12552 2834 12608
rect 2502 9832 2558 9888
rect 2318 9424 2374 9480
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 3606 16360 3662 16416
rect 3698 16088 3754 16144
rect 3698 15680 3754 15736
rect 4342 16360 4398 16416
rect 3606 14184 3662 14240
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 2870 11328 2926 11384
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 3974 14320 4030 14376
rect 4526 15020 4582 15056
rect 4526 15000 4528 15020
rect 4528 15000 4580 15020
rect 4580 15000 4582 15020
rect 4618 14764 4620 14784
rect 4620 14764 4672 14784
rect 4672 14764 4674 14784
rect 4618 14728 4674 14764
rect 3882 13368 3938 13424
rect 3790 13232 3846 13288
rect 3698 12824 3754 12880
rect 3606 11872 3662 11928
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 4802 15952 4858 16008
rect 4710 13504 4766 13560
rect 4710 13368 4766 13424
rect 4710 12960 4766 13016
rect 5446 16532 5448 16552
rect 5448 16532 5500 16552
rect 5500 16532 5502 16552
rect 5446 16496 5502 16532
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 5538 15036 5540 15056
rect 5540 15036 5592 15056
rect 5592 15036 5594 15056
rect 5538 15000 5594 15036
rect 4710 12708 4766 12744
rect 5354 14864 5410 14920
rect 5262 14340 5318 14376
rect 5262 14320 5264 14340
rect 5264 14320 5316 14340
rect 5316 14320 5318 14340
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 4710 12688 4712 12708
rect 4712 12688 4764 12708
rect 4764 12688 4766 12708
rect 4342 12144 4398 12200
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 2962 9968 3018 10024
rect 2870 9424 2926 9480
rect 3422 9424 3478 9480
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 3514 8880 3570 8936
rect 2962 8064 3018 8120
rect 2778 6840 2834 6896
rect 1582 5208 1638 5264
rect 2870 6432 2926 6488
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 2962 6024 3018 6080
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3974 10512 4030 10568
rect 3882 9968 3938 10024
rect 3698 9152 3754 9208
rect 4434 11464 4490 11520
rect 4158 9988 4214 10024
rect 4158 9968 4160 9988
rect 4160 9968 4212 9988
rect 4212 9968 4214 9988
rect 4066 9580 4122 9616
rect 4066 9560 4068 9580
rect 4068 9560 4120 9580
rect 4120 9560 4122 9580
rect 4250 9424 4306 9480
rect 4434 10648 4490 10704
rect 4526 10376 4582 10432
rect 4158 9288 4214 9344
rect 4066 8472 4122 8528
rect 4342 9152 4398 9208
rect 4250 8744 4306 8800
rect 4066 7656 4122 7712
rect 3974 7248 4030 7304
rect 4986 12688 5042 12744
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 5262 12280 5318 12336
rect 4986 12164 5042 12200
rect 4986 12144 4988 12164
rect 4988 12144 5040 12164
rect 5040 12144 5042 12164
rect 5998 16632 6054 16688
rect 5998 15272 6054 15328
rect 5906 13776 5962 13832
rect 6182 14456 6238 14512
rect 6274 14320 6330 14376
rect 5814 12960 5870 13016
rect 3974 5652 3976 5672
rect 3976 5652 4028 5672
rect 4028 5652 4030 5672
rect 3974 5616 4030 5652
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 5078 11736 5134 11792
rect 5354 11620 5410 11656
rect 5354 11600 5356 11620
rect 5356 11600 5408 11620
rect 5408 11600 5410 11620
rect 5170 10956 5172 10976
rect 5172 10956 5224 10976
rect 5224 10956 5226 10976
rect 5170 10920 5226 10956
rect 5170 10376 5226 10432
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 5538 10668 5594 10704
rect 5538 10648 5540 10668
rect 5540 10648 5592 10668
rect 5592 10648 5594 10668
rect 5446 9988 5502 10024
rect 5446 9968 5448 9988
rect 5448 9968 5500 9988
rect 5500 9968 5502 9988
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 5630 9560 5686 9616
rect 5262 9288 5318 9344
rect 5538 9172 5594 9208
rect 5538 9152 5540 9172
rect 5540 9152 5592 9172
rect 5592 9152 5594 9172
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 5262 8084 5318 8120
rect 5262 8064 5264 8084
rect 5264 8064 5316 8084
rect 5316 8064 5318 8084
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 5998 12960 6054 13016
rect 5814 7404 5870 7440
rect 5814 7384 5816 7404
rect 5816 7384 5868 7404
rect 5868 7384 5870 7404
rect 6458 13812 6460 13832
rect 6460 13812 6512 13832
rect 6512 13812 6514 13832
rect 6458 13776 6514 13812
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 6182 9016 6238 9072
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 7194 16224 7250 16280
rect 7194 13640 7250 13696
rect 7010 11464 7066 11520
rect 6642 9424 6698 9480
rect 6826 9172 6882 9208
rect 6826 9152 6828 9172
rect 6828 9152 6880 9172
rect 6880 9152 6882 9172
rect 7838 15952 7894 16008
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 7470 15000 7526 15056
rect 7746 15444 7748 15464
rect 7748 15444 7800 15464
rect 7800 15444 7802 15464
rect 7746 15408 7802 15444
rect 7838 15136 7894 15192
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 7654 13368 7710 13424
rect 7654 12724 7656 12744
rect 7656 12724 7708 12744
rect 7708 12724 7710 12744
rect 7654 12688 7710 12724
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 7194 11056 7250 11112
rect 8206 16224 8262 16280
rect 8114 15816 8170 15872
rect 8114 15136 8170 15192
rect 8022 14456 8078 14512
rect 8298 15816 8354 15872
rect 8298 14864 8354 14920
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 8666 15952 8722 16008
rect 8206 13232 8262 13288
rect 8482 13812 8484 13832
rect 8484 13812 8536 13832
rect 8536 13812 8538 13832
rect 8482 13776 8538 13812
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 9310 15408 9366 15464
rect 9218 15272 9274 15328
rect 9126 12316 9128 12336
rect 9128 12316 9180 12336
rect 9180 12316 9182 12336
rect 9126 12280 9182 12316
rect 8666 10668 8722 10704
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 9402 13388 9458 13424
rect 9402 13368 9404 13388
rect 9404 13368 9456 13388
rect 9456 13368 9458 13388
rect 9862 13232 9918 13288
rect 9310 12824 9366 12880
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 9678 12824 9734 12880
rect 10138 12416 10194 12472
rect 10046 12280 10102 12336
rect 10230 12144 10286 12200
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 8666 10648 8668 10668
rect 8668 10648 8720 10668
rect 8720 10648 8722 10668
rect 9126 10260 9182 10296
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 10506 15136 10562 15192
rect 10506 14884 10562 14920
rect 10506 14864 10508 14884
rect 10508 14864 10560 14884
rect 10560 14864 10562 14884
rect 10690 15444 10692 15464
rect 10692 15444 10744 15464
rect 10744 15444 10746 15464
rect 10690 15408 10746 15444
rect 10690 15308 10692 15328
rect 10692 15308 10744 15328
rect 10744 15308 10746 15328
rect 10690 15272 10746 15308
rect 10782 15000 10838 15056
rect 10414 13368 10470 13424
rect 10506 12416 10562 12472
rect 9126 10240 9128 10260
rect 9128 10240 9180 10260
rect 9180 10240 9182 10260
rect 8666 9580 8722 9616
rect 8666 9560 8668 9580
rect 8668 9560 8720 9580
rect 8720 9560 8722 9580
rect 9126 9580 9182 9616
rect 9126 9560 9128 9580
rect 9128 9560 9180 9580
rect 9180 9560 9182 9580
rect 8114 9424 8170 9480
rect 7194 8492 7250 8528
rect 7194 8472 7196 8492
rect 7196 8472 7248 8492
rect 7248 8472 7250 8492
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 11150 11736 11206 11792
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 12438 15136 12494 15192
rect 12162 14864 12218 14920
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 13082 15952 13138 16008
rect 12990 15272 13046 15328
rect 13358 15544 13414 15600
rect 12898 13776 12954 13832
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 11702 11756 11758 11792
rect 11702 11736 11704 11756
rect 11704 11736 11756 11756
rect 11756 11736 11758 11756
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 11058 11228 11060 11248
rect 11060 11228 11112 11248
rect 11112 11228 11114 11248
rect 11058 11192 11114 11228
rect 13542 15000 13598 15056
rect 13818 14320 13874 14376
rect 13910 13504 13966 13560
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 14370 15544 14426 15600
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 14922 15988 14924 16008
rect 14924 15988 14976 16008
rect 14976 15988 14978 16008
rect 14922 15952 14978 15988
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 14370 13912 14426 13968
rect 13726 11756 13782 11792
rect 13726 11736 13728 11756
rect 13728 11736 13780 11756
rect 13780 11736 13782 11756
rect 14554 13676 14556 13696
rect 14556 13676 14608 13696
rect 14608 13676 14610 13696
rect 14554 13640 14610 13676
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 14462 11328 14518 11384
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 15014 15444 15016 15464
rect 15016 15444 15068 15464
rect 15068 15444 15070 15464
rect 15014 15408 15070 15444
rect 16026 18944 16082 19000
rect 15290 16516 15346 16552
rect 15290 16496 15292 16516
rect 15292 16496 15344 16516
rect 15344 16496 15346 16516
rect 15198 14048 15254 14104
rect 15658 15544 15714 15600
rect 15290 13640 15346 13696
rect 15474 13640 15530 13696
rect 15382 12960 15438 13016
rect 15474 12824 15530 12880
rect 15474 12552 15530 12608
rect 15842 17040 15898 17096
rect 15658 13368 15714 13424
rect 15842 14184 15898 14240
rect 15658 13232 15714 13288
rect 15750 13096 15806 13152
rect 16394 17720 16450 17776
rect 16026 15000 16082 15056
rect 16026 14864 16082 14920
rect 16026 13368 16082 13424
rect 16210 15952 16266 16008
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 16394 15000 16450 15056
rect 16210 14728 16266 14784
rect 16210 14220 16212 14240
rect 16212 14220 16264 14240
rect 16264 14220 16266 14240
rect 16210 14184 16266 14220
rect 16210 13640 16266 13696
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 16486 14320 16542 14376
rect 17130 15408 17186 15464
rect 17038 14320 17094 14376
rect 16486 13776 16542 13832
rect 16670 13776 16726 13832
rect 16946 14048 17002 14104
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 16946 13776 17002 13832
rect 16946 12824 17002 12880
rect 16302 12708 16358 12744
rect 16302 12688 16304 12708
rect 16304 12688 16356 12708
rect 16356 12688 16358 12708
rect 16210 12416 16266 12472
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 17498 11620 17554 11656
rect 17498 11600 17500 11620
rect 17500 11600 17552 11620
rect 17552 11600 17554 11620
rect 17682 14456 17738 14512
rect 19062 18128 19118 18184
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 18602 16088 18658 16144
rect 17958 13504 18014 13560
rect 18234 13504 18290 13560
rect 17958 11756 18014 11792
rect 17958 11736 17960 11756
rect 17960 11736 18012 11756
rect 18012 11736 18014 11756
rect 17682 10648 17738 10704
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 18326 11192 18382 11248
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 18510 11736 18566 11792
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 18326 10376 18382 10432
rect 18326 9968 18382 10024
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 18326 9172 18382 9208
rect 18326 9152 18328 9172
rect 18328 9152 18380 9172
rect 18380 9152 18382 9172
rect 19154 8744 19210 8800
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 18326 7948 18382 7984
rect 18326 7928 18328 7948
rect 18328 7928 18380 7948
rect 18380 7928 18382 7948
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 18326 7404 18382 7440
rect 18326 7384 18328 7404
rect 18328 7384 18380 7404
rect 18380 7384 18382 7404
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 18326 6740 18328 6760
rect 18328 6740 18380 6760
rect 18380 6740 18382 6760
rect 18326 6704 18382 6740
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 18326 6316 18382 6352
rect 18326 6296 18328 6316
rect 18328 6296 18380 6316
rect 18380 6296 18382 6316
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 18326 5652 18328 5672
rect 18328 5652 18380 5672
rect 18380 5652 18382 5672
rect 18326 5616 18382 5652
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 18326 5092 18382 5128
rect 18326 5072 18328 5092
rect 18328 5072 18380 5092
rect 18380 5072 18382 5092
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 1674 4428 1676 4448
rect 1676 4428 1728 4448
rect 1728 4428 1730 4448
rect 1674 4392 1730 4428
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 19154 4256 19210 4312
rect 1582 3984 1638 4040
rect 18326 3884 18328 3904
rect 18328 3884 18380 3904
rect 18380 3884 18382 3904
rect 18326 3848 18382 3884
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 1582 3168 1638 3224
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 18326 3032 18382 3088
rect 1582 2760 1638 2816
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 18326 2624 18382 2680
rect 2226 1944 2282 2000
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 2870 1536 2926 1592
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
rect 18326 1808 18382 1864
rect 17682 1400 17738 1456
<< metal3 >>
rect 16021 19002 16087 19005
rect 19200 19002 20000 19032
rect 16021 19000 20000 19002
rect 16021 18944 16026 19000
rect 16082 18944 20000 19000
rect 16021 18942 20000 18944
rect 16021 18939 16087 18942
rect 19200 18912 20000 18942
rect 381 18594 447 18597
rect 7230 18594 7236 18596
rect 381 18592 7236 18594
rect 381 18536 386 18592
rect 442 18536 7236 18592
rect 381 18534 7236 18536
rect 381 18531 447 18534
rect 7230 18532 7236 18534
rect 7300 18532 7306 18596
rect 13670 18532 13676 18596
rect 13740 18594 13746 18596
rect 19200 18594 20000 18624
rect 13740 18534 20000 18594
rect 13740 18532 13746 18534
rect 19200 18504 20000 18534
rect 0 18322 800 18352
rect 6126 18322 6132 18324
rect 0 18262 6132 18322
rect 0 18232 800 18262
rect 6126 18260 6132 18262
rect 6196 18260 6202 18324
rect 19057 18186 19123 18189
rect 19200 18186 20000 18216
rect 19057 18184 20000 18186
rect 19057 18128 19062 18184
rect 19118 18128 20000 18184
rect 19057 18126 20000 18128
rect 19057 18123 19123 18126
rect 19200 18096 20000 18126
rect 0 17914 800 17944
rect 9254 17914 9260 17916
rect 0 17854 9260 17914
rect 0 17824 800 17854
rect 9254 17852 9260 17854
rect 9324 17852 9330 17916
rect 16389 17778 16455 17781
rect 19200 17778 20000 17808
rect 16389 17776 20000 17778
rect 16389 17720 16394 17776
rect 16450 17720 20000 17776
rect 16389 17718 20000 17720
rect 16389 17715 16455 17718
rect 19200 17688 20000 17718
rect 0 17506 800 17536
rect 0 17446 2790 17506
rect 0 17416 800 17446
rect 2730 17234 2790 17446
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 19200 17370 20000 17400
rect 19152 17280 20000 17370
rect 7414 17234 7420 17236
rect 2730 17174 7420 17234
rect 7414 17172 7420 17174
rect 7484 17172 7490 17236
rect 14774 17172 14780 17236
rect 14844 17234 14850 17236
rect 19152 17234 19212 17280
rect 14844 17174 19212 17234
rect 14844 17172 14850 17174
rect 0 17098 800 17128
rect 2037 17098 2103 17101
rect 11462 17098 11468 17100
rect 0 17096 2103 17098
rect 0 17040 2042 17096
rect 2098 17040 2103 17096
rect 0 17038 2103 17040
rect 0 17008 800 17038
rect 2037 17035 2103 17038
rect 5812 17038 11468 17098
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 0 16690 800 16720
rect 5812 16690 5872 17038
rect 11462 17036 11468 17038
rect 11532 17036 11538 17100
rect 15837 17098 15903 17101
rect 15837 17096 17050 17098
rect 15837 17040 15842 17096
rect 15898 17040 17050 17096
rect 15837 17038 17050 17040
rect 15837 17035 15903 17038
rect 16990 16962 17050 17038
rect 19200 16962 20000 16992
rect 16990 16902 20000 16962
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 19200 16872 20000 16902
rect 16482 16831 16798 16832
rect 0 16630 5872 16690
rect 5993 16690 6059 16693
rect 10358 16690 10364 16692
rect 5993 16688 10364 16690
rect 5993 16632 5998 16688
rect 6054 16632 10364 16688
rect 5993 16630 10364 16632
rect 0 16600 800 16630
rect 5993 16627 6059 16630
rect 10358 16628 10364 16630
rect 10428 16628 10434 16692
rect 5441 16554 5507 16557
rect 9070 16554 9076 16556
rect 5441 16552 9076 16554
rect 5441 16496 5446 16552
rect 5502 16496 9076 16552
rect 5441 16494 9076 16496
rect 5441 16491 5507 16494
rect 9070 16492 9076 16494
rect 9140 16492 9146 16556
rect 15285 16554 15351 16557
rect 19200 16554 20000 16584
rect 15285 16552 20000 16554
rect 15285 16496 15290 16552
rect 15346 16496 20000 16552
rect 15285 16494 20000 16496
rect 15285 16491 15351 16494
rect 19200 16464 20000 16494
rect 3601 16418 3667 16421
rect 4337 16418 4403 16421
rect 3601 16416 4403 16418
rect 3601 16360 3606 16416
rect 3662 16360 4342 16416
rect 4398 16360 4403 16416
rect 3601 16358 4403 16360
rect 3601 16355 3667 16358
rect 4337 16355 4403 16358
rect 5384 16352 5700 16353
rect 0 16282 800 16312
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 4286 16282 4292 16284
rect 0 16222 4292 16282
rect 0 16192 800 16222
rect 4286 16220 4292 16222
rect 4356 16220 4362 16284
rect 7189 16282 7255 16285
rect 8201 16282 8267 16285
rect 7189 16280 8267 16282
rect 7189 16224 7194 16280
rect 7250 16224 8206 16280
rect 8262 16224 8267 16280
rect 7189 16222 8267 16224
rect 7189 16219 7255 16222
rect 8201 16219 8267 16222
rect 3693 16146 3759 16149
rect 8150 16146 8156 16148
rect 3693 16144 8156 16146
rect 3693 16088 3698 16144
rect 3754 16088 8156 16144
rect 3693 16086 8156 16088
rect 3693 16083 3759 16086
rect 8150 16084 8156 16086
rect 8220 16084 8226 16148
rect 18597 16146 18663 16149
rect 19200 16146 20000 16176
rect 18597 16144 20000 16146
rect 18597 16088 18602 16144
rect 18658 16088 20000 16144
rect 18597 16086 20000 16088
rect 18597 16083 18663 16086
rect 19200 16056 20000 16086
rect 4797 16010 4863 16013
rect 5206 16010 5212 16012
rect 4797 16008 5212 16010
rect 4797 15952 4802 16008
rect 4858 15952 5212 16008
rect 4797 15950 5212 15952
rect 4797 15947 4863 15950
rect 5206 15948 5212 15950
rect 5276 15948 5282 16012
rect 7833 16010 7899 16013
rect 8661 16010 8727 16013
rect 7833 16008 8727 16010
rect 7833 15952 7838 16008
rect 7894 15952 8666 16008
rect 8722 15952 8727 16008
rect 7833 15950 8727 15952
rect 7833 15947 7899 15950
rect 8661 15947 8727 15950
rect 13077 16010 13143 16013
rect 14917 16010 14983 16013
rect 16205 16010 16271 16013
rect 13077 16008 16271 16010
rect 13077 15952 13082 16008
rect 13138 15952 14922 16008
rect 14978 15952 16210 16008
rect 16266 15952 16271 16008
rect 13077 15950 16271 15952
rect 13077 15947 13143 15950
rect 14917 15947 14983 15950
rect 16205 15947 16271 15950
rect 0 15874 800 15904
rect 8109 15874 8175 15877
rect 8293 15874 8359 15877
rect 0 15814 2790 15874
rect 0 15784 800 15814
rect 2730 15602 2790 15814
rect 8109 15872 8359 15874
rect 8109 15816 8114 15872
rect 8170 15816 8298 15872
rect 8354 15816 8359 15872
rect 8109 15814 8359 15816
rect 8109 15811 8175 15814
rect 8293 15811 8359 15814
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 3693 15738 3759 15741
rect 19200 15738 20000 15768
rect 3693 15736 7298 15738
rect 3693 15680 3698 15736
rect 3754 15680 7298 15736
rect 3693 15678 7298 15680
rect 3693 15675 3759 15678
rect 7046 15602 7052 15604
rect 2730 15542 7052 15602
rect 7046 15540 7052 15542
rect 7116 15540 7122 15604
rect 7238 15602 7298 15678
rect 16990 15678 20000 15738
rect 9622 15602 9628 15604
rect 7238 15542 9628 15602
rect 9622 15540 9628 15542
rect 9692 15540 9698 15604
rect 13353 15602 13419 15605
rect 14365 15602 14431 15605
rect 13353 15600 14431 15602
rect 13353 15544 13358 15600
rect 13414 15544 14370 15600
rect 14426 15544 14431 15600
rect 13353 15542 14431 15544
rect 13353 15539 13419 15542
rect 14365 15539 14431 15542
rect 15653 15602 15719 15605
rect 16990 15602 17050 15678
rect 19200 15648 20000 15678
rect 15653 15600 17050 15602
rect 15653 15544 15658 15600
rect 15714 15544 17050 15600
rect 15653 15542 17050 15544
rect 15653 15539 15719 15542
rect 0 15466 800 15496
rect 2957 15466 3023 15469
rect 0 15464 3023 15466
rect 0 15408 2962 15464
rect 3018 15408 3023 15464
rect 0 15406 3023 15408
rect 0 15376 800 15406
rect 2957 15403 3023 15406
rect 7741 15466 7807 15469
rect 9305 15466 9371 15469
rect 7741 15464 9371 15466
rect 7741 15408 7746 15464
rect 7802 15408 9310 15464
rect 9366 15408 9371 15464
rect 7741 15406 9371 15408
rect 7741 15403 7807 15406
rect 9305 15403 9371 15406
rect 10542 15404 10548 15468
rect 10612 15466 10618 15468
rect 10685 15466 10751 15469
rect 10612 15464 10751 15466
rect 10612 15408 10690 15464
rect 10746 15408 10751 15464
rect 10612 15406 10751 15408
rect 10612 15404 10618 15406
rect 10685 15403 10751 15406
rect 15009 15466 15075 15469
rect 17125 15466 17191 15469
rect 15009 15464 17191 15466
rect 15009 15408 15014 15464
rect 15070 15408 17130 15464
rect 17186 15408 17191 15464
rect 15009 15406 17191 15408
rect 15009 15403 15075 15406
rect 17125 15403 17191 15406
rect 17358 15406 19212 15466
rect 5993 15330 6059 15333
rect 9213 15330 9279 15333
rect 5993 15328 9279 15330
rect 5993 15272 5998 15328
rect 6054 15272 9218 15328
rect 9274 15272 9279 15328
rect 5993 15270 9279 15272
rect 5993 15267 6059 15270
rect 9213 15267 9279 15270
rect 10685 15330 10751 15333
rect 12985 15330 13051 15333
rect 10685 15328 13051 15330
rect 10685 15272 10690 15328
rect 10746 15272 12990 15328
rect 13046 15272 13051 15328
rect 10685 15270 13051 15272
rect 10685 15267 10751 15270
rect 12985 15267 13051 15270
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 7833 15194 7899 15197
rect 8109 15194 8175 15197
rect 7833 15192 8175 15194
rect 7833 15136 7838 15192
rect 7894 15136 8114 15192
rect 8170 15136 8175 15192
rect 7833 15134 8175 15136
rect 7833 15131 7899 15134
rect 8109 15131 8175 15134
rect 10501 15194 10567 15197
rect 12433 15194 12499 15197
rect 17358 15194 17418 15406
rect 19152 15360 19212 15406
rect 19152 15270 20000 15360
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 19200 15240 20000 15270
rect 18701 15199 19017 15200
rect 10501 15192 12499 15194
rect 10501 15136 10506 15192
rect 10562 15136 12438 15192
rect 12494 15136 12499 15192
rect 10501 15134 12499 15136
rect 10501 15131 10567 15134
rect 12433 15131 12499 15134
rect 14782 15134 17418 15194
rect 0 15058 800 15088
rect 2865 15058 2931 15061
rect 0 15056 2931 15058
rect 0 15000 2870 15056
rect 2926 15000 2931 15056
rect 0 14998 2931 15000
rect 0 14968 800 14998
rect 2865 14995 2931 14998
rect 4521 15058 4587 15061
rect 5533 15058 5599 15061
rect 4521 15056 5599 15058
rect 4521 15000 4526 15056
rect 4582 15000 5538 15056
rect 5594 15000 5599 15056
rect 4521 14998 5599 15000
rect 4521 14995 4587 14998
rect 5533 14995 5599 14998
rect 7465 15058 7531 15061
rect 10777 15058 10843 15061
rect 7465 15056 10843 15058
rect 7465 15000 7470 15056
rect 7526 15000 10782 15056
rect 10838 15000 10843 15056
rect 7465 14998 10843 15000
rect 7465 14995 7531 14998
rect 10777 14995 10843 14998
rect 13537 15058 13603 15061
rect 14782 15058 14842 15134
rect 13537 15056 14842 15058
rect 13537 15000 13542 15056
rect 13598 15000 14842 15056
rect 13537 14998 14842 15000
rect 13537 14995 13603 14998
rect 15878 14996 15884 15060
rect 15948 15058 15954 15060
rect 16021 15058 16087 15061
rect 15948 15056 16087 15058
rect 15948 15000 16026 15056
rect 16082 15000 16087 15056
rect 15948 14998 16087 15000
rect 15948 14996 15954 14998
rect 16021 14995 16087 14998
rect 16246 14996 16252 15060
rect 16316 15058 16322 15060
rect 16389 15058 16455 15061
rect 16316 15056 16455 15058
rect 16316 15000 16394 15056
rect 16450 15000 16455 15056
rect 16316 14998 16455 15000
rect 16316 14996 16322 14998
rect 16389 14995 16455 14998
rect 5349 14922 5415 14925
rect 8293 14922 8359 14925
rect 5349 14920 8359 14922
rect 5349 14864 5354 14920
rect 5410 14864 8298 14920
rect 8354 14864 8359 14920
rect 5349 14862 8359 14864
rect 5349 14859 5415 14862
rect 8293 14859 8359 14862
rect 10501 14922 10567 14925
rect 12157 14922 12223 14925
rect 10501 14920 12223 14922
rect 10501 14864 10506 14920
rect 10562 14864 12162 14920
rect 12218 14864 12223 14920
rect 10501 14862 12223 14864
rect 10501 14859 10567 14862
rect 12157 14859 12223 14862
rect 16021 14922 16087 14925
rect 19200 14922 20000 14952
rect 16021 14920 20000 14922
rect 16021 14864 16026 14920
rect 16082 14864 20000 14920
rect 16021 14862 20000 14864
rect 16021 14859 16087 14862
rect 19200 14832 20000 14862
rect 4470 14724 4476 14788
rect 4540 14786 4546 14788
rect 4613 14786 4679 14789
rect 4540 14784 4679 14786
rect 4540 14728 4618 14784
rect 4674 14728 4679 14784
rect 4540 14726 4679 14728
rect 4540 14724 4546 14726
rect 4613 14723 4679 14726
rect 16062 14724 16068 14788
rect 16132 14786 16138 14788
rect 16205 14786 16271 14789
rect 16132 14784 16271 14786
rect 16132 14728 16210 14784
rect 16266 14728 16271 14784
rect 16132 14726 16271 14728
rect 16132 14724 16138 14726
rect 16205 14723 16271 14726
rect 3165 14720 3481 14721
rect 0 14650 800 14680
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 2998 14650 3004 14652
rect 0 14590 3004 14650
rect 0 14560 800 14590
rect 2998 14588 3004 14590
rect 3068 14588 3074 14652
rect 6177 14514 6243 14517
rect 8017 14514 8083 14517
rect 6177 14512 8083 14514
rect 6177 14456 6182 14512
rect 6238 14456 8022 14512
rect 8078 14456 8083 14512
rect 6177 14454 8083 14456
rect 6177 14451 6243 14454
rect 8017 14451 8083 14454
rect 17677 14514 17743 14517
rect 19200 14514 20000 14544
rect 17677 14512 20000 14514
rect 17677 14456 17682 14512
rect 17738 14456 20000 14512
rect 17677 14454 20000 14456
rect 17677 14451 17743 14454
rect 19200 14424 20000 14454
rect 3969 14378 4035 14381
rect 5257 14378 5323 14381
rect 6269 14378 6335 14381
rect 3969 14376 6335 14378
rect 3969 14320 3974 14376
rect 4030 14320 5262 14376
rect 5318 14320 6274 14376
rect 6330 14320 6335 14376
rect 3969 14318 6335 14320
rect 3969 14315 4035 14318
rect 5257 14315 5323 14318
rect 6269 14315 6335 14318
rect 13813 14378 13879 14381
rect 16481 14378 16547 14381
rect 17033 14378 17099 14381
rect 17902 14378 17908 14380
rect 13813 14376 17908 14378
rect 13813 14320 13818 14376
rect 13874 14320 16486 14376
rect 16542 14320 17038 14376
rect 17094 14320 17908 14376
rect 13813 14318 17908 14320
rect 13813 14315 13879 14318
rect 16481 14315 16547 14318
rect 17033 14315 17099 14318
rect 17902 14316 17908 14318
rect 17972 14316 17978 14380
rect 0 14242 800 14272
rect 3601 14242 3667 14245
rect 0 14240 3667 14242
rect 0 14184 3606 14240
rect 3662 14184 3667 14240
rect 0 14182 3667 14184
rect 0 14152 800 14182
rect 3601 14179 3667 14182
rect 15837 14242 15903 14245
rect 16205 14242 16271 14245
rect 15837 14240 16271 14242
rect 15837 14184 15842 14240
rect 15898 14184 16210 14240
rect 16266 14184 16271 14240
rect 15837 14182 16271 14184
rect 15837 14179 15903 14182
rect 16205 14179 16271 14182
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 15193 14106 15259 14109
rect 16941 14106 17007 14109
rect 19200 14106 20000 14136
rect 15193 14104 17007 14106
rect 15193 14048 15198 14104
rect 15254 14048 16946 14104
rect 17002 14048 17007 14104
rect 15193 14046 17007 14048
rect 15193 14043 15259 14046
rect 16941 14043 17007 14046
rect 19152 14016 20000 14106
rect 2589 13970 2655 13973
rect 4102 13970 4108 13972
rect 2589 13968 4108 13970
rect 2589 13912 2594 13968
rect 2650 13912 4108 13968
rect 2589 13910 4108 13912
rect 2589 13907 2655 13910
rect 4102 13908 4108 13910
rect 4172 13908 4178 13972
rect 14365 13970 14431 13973
rect 19152 13970 19212 14016
rect 14365 13968 19212 13970
rect 14365 13912 14370 13968
rect 14426 13912 19212 13968
rect 14365 13910 19212 13912
rect 14365 13907 14431 13910
rect 0 13834 800 13864
rect 5901 13834 5967 13837
rect 6453 13834 6519 13837
rect 8477 13834 8543 13837
rect 0 13774 5826 13834
rect 0 13744 800 13774
rect 5766 13698 5826 13774
rect 5901 13832 8543 13834
rect 5901 13776 5906 13832
rect 5962 13776 6458 13832
rect 6514 13776 8482 13832
rect 8538 13776 8543 13832
rect 5901 13774 8543 13776
rect 5901 13771 5967 13774
rect 6453 13771 6519 13774
rect 8477 13771 8543 13774
rect 12893 13834 12959 13837
rect 16481 13834 16547 13837
rect 12893 13832 16547 13834
rect 12893 13776 12898 13832
rect 12954 13776 16486 13832
rect 16542 13776 16547 13832
rect 12893 13774 16547 13776
rect 12893 13771 12959 13774
rect 16481 13771 16547 13774
rect 16665 13834 16731 13837
rect 16941 13834 17007 13837
rect 16665 13832 17007 13834
rect 16665 13776 16670 13832
rect 16726 13776 16946 13832
rect 17002 13776 17007 13832
rect 16665 13774 17007 13776
rect 16665 13771 16731 13774
rect 16941 13771 17007 13774
rect 7189 13698 7255 13701
rect 5766 13696 7255 13698
rect 5766 13640 7194 13696
rect 7250 13640 7255 13696
rect 5766 13638 7255 13640
rect 7189 13635 7255 13638
rect 14549 13698 14615 13701
rect 15285 13698 15351 13701
rect 14549 13696 15351 13698
rect 14549 13640 14554 13696
rect 14610 13640 15290 13696
rect 15346 13640 15351 13696
rect 14549 13638 15351 13640
rect 14549 13635 14615 13638
rect 15285 13635 15351 13638
rect 15469 13698 15535 13701
rect 16205 13698 16271 13701
rect 19200 13698 20000 13728
rect 15469 13696 16271 13698
rect 15469 13640 15474 13696
rect 15530 13640 16210 13696
rect 16266 13640 16271 13696
rect 15469 13638 16271 13640
rect 15469 13635 15535 13638
rect 16205 13635 16271 13638
rect 17726 13638 20000 13698
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 4705 13562 4771 13565
rect 6678 13562 6684 13564
rect 4705 13560 6684 13562
rect 4705 13504 4710 13560
rect 4766 13504 6684 13560
rect 4705 13502 6684 13504
rect 4705 13499 4771 13502
rect 6678 13500 6684 13502
rect 6748 13500 6754 13564
rect 13905 13562 13971 13565
rect 15472 13562 15532 13635
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 13905 13560 15532 13562
rect 13905 13504 13910 13560
rect 13966 13504 15532 13560
rect 13905 13502 15532 13504
rect 13905 13499 13971 13502
rect 0 13426 800 13456
rect 3877 13426 3943 13429
rect 0 13424 3943 13426
rect 0 13368 3882 13424
rect 3938 13368 3943 13424
rect 0 13366 3943 13368
rect 0 13336 800 13366
rect 3877 13363 3943 13366
rect 4705 13426 4771 13429
rect 7649 13426 7715 13429
rect 4705 13424 7715 13426
rect 4705 13368 4710 13424
rect 4766 13368 7654 13424
rect 7710 13368 7715 13424
rect 4705 13366 7715 13368
rect 4705 13363 4771 13366
rect 7649 13363 7715 13366
rect 9397 13426 9463 13429
rect 10409 13426 10475 13429
rect 15653 13426 15719 13429
rect 9397 13424 10475 13426
rect 9397 13368 9402 13424
rect 9458 13368 10414 13424
rect 10470 13368 10475 13424
rect 9397 13366 10475 13368
rect 9397 13363 9463 13366
rect 10409 13363 10475 13366
rect 15518 13424 15719 13426
rect 15518 13368 15658 13424
rect 15714 13368 15719 13424
rect 15518 13366 15719 13368
rect 3785 13290 3851 13293
rect 8201 13290 8267 13293
rect 3785 13288 8267 13290
rect 3785 13232 3790 13288
rect 3846 13232 8206 13288
rect 8262 13232 8267 13288
rect 3785 13230 8267 13232
rect 3785 13227 3851 13230
rect 8201 13227 8267 13230
rect 9857 13290 9923 13293
rect 9857 13288 12956 13290
rect 9857 13232 9862 13288
rect 9918 13232 12956 13288
rect 9857 13230 12956 13232
rect 9857 13227 9923 13230
rect 5384 13088 5700 13089
rect 0 13018 800 13048
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 4705 13018 4771 13021
rect 0 13016 4771 13018
rect 0 12960 4710 13016
rect 4766 12960 4771 13016
rect 0 12958 4771 12960
rect 0 12928 800 12958
rect 4705 12955 4771 12958
rect 5809 13018 5875 13021
rect 5993 13018 6059 13021
rect 5809 13016 6059 13018
rect 5809 12960 5814 13016
rect 5870 12960 5998 13016
rect 6054 12960 6059 13016
rect 5809 12958 6059 12960
rect 5809 12955 5875 12958
rect 5993 12955 6059 12958
rect 3693 12882 3759 12885
rect 9305 12882 9371 12885
rect 3693 12880 9371 12882
rect 3693 12824 3698 12880
rect 3754 12824 9310 12880
rect 9366 12824 9371 12880
rect 3693 12822 9371 12824
rect 3693 12819 3759 12822
rect 9305 12819 9371 12822
rect 9673 12882 9739 12885
rect 10542 12882 10548 12884
rect 9673 12880 10548 12882
rect 9673 12824 9678 12880
rect 9734 12824 10548 12880
rect 9673 12822 10548 12824
rect 9673 12819 9739 12822
rect 10542 12820 10548 12822
rect 10612 12820 10618 12884
rect 12896 12882 12956 13230
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 15377 13018 15443 13021
rect 15518 13018 15578 13366
rect 15653 13363 15719 13366
rect 16021 13426 16087 13429
rect 17726 13426 17786 13638
rect 19200 13608 20000 13638
rect 17953 13562 18019 13565
rect 18229 13562 18295 13565
rect 17953 13560 18295 13562
rect 17953 13504 17958 13560
rect 18014 13504 18234 13560
rect 18290 13504 18295 13560
rect 17953 13502 18295 13504
rect 17953 13499 18019 13502
rect 18229 13499 18295 13502
rect 16021 13424 17786 13426
rect 16021 13368 16026 13424
rect 16082 13368 17786 13424
rect 16021 13366 17786 13368
rect 16021 13363 16087 13366
rect 15653 13290 15719 13293
rect 19200 13290 20000 13320
rect 15653 13288 20000 13290
rect 15653 13232 15658 13288
rect 15714 13232 20000 13288
rect 15653 13230 20000 13232
rect 15653 13227 15719 13230
rect 19200 13200 20000 13230
rect 15745 13154 15811 13157
rect 15878 13154 15884 13156
rect 15745 13152 15884 13154
rect 15745 13096 15750 13152
rect 15806 13096 15884 13152
rect 15745 13094 15884 13096
rect 15745 13091 15811 13094
rect 15878 13092 15884 13094
rect 15948 13092 15954 13156
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 15377 13016 15578 13018
rect 15377 12960 15382 13016
rect 15438 12960 15578 13016
rect 15377 12958 15578 12960
rect 15377 12955 15443 12958
rect 15469 12882 15535 12885
rect 12896 12880 15535 12882
rect 12896 12824 15474 12880
rect 15530 12824 15535 12880
rect 12896 12822 15535 12824
rect 15469 12819 15535 12822
rect 16941 12882 17007 12885
rect 19200 12882 20000 12912
rect 16941 12880 20000 12882
rect 16941 12824 16946 12880
rect 17002 12824 20000 12880
rect 16941 12822 20000 12824
rect 16941 12819 17007 12822
rect 19200 12792 20000 12822
rect 2681 12746 2747 12749
rect 4705 12746 4771 12749
rect 2681 12744 4771 12746
rect 2681 12688 2686 12744
rect 2742 12688 4710 12744
rect 4766 12688 4771 12744
rect 2681 12686 4771 12688
rect 2681 12683 2747 12686
rect 4705 12683 4771 12686
rect 4981 12746 5047 12749
rect 7649 12746 7715 12749
rect 4981 12744 7715 12746
rect 4981 12688 4986 12744
rect 5042 12688 7654 12744
rect 7710 12688 7715 12744
rect 4981 12686 7715 12688
rect 4981 12683 5047 12686
rect 7649 12683 7715 12686
rect 16297 12746 16363 12749
rect 16297 12744 17832 12746
rect 16297 12688 16302 12744
rect 16358 12688 17832 12744
rect 16297 12686 17832 12688
rect 16297 12683 16363 12686
rect 0 12610 800 12640
rect 2773 12610 2839 12613
rect 0 12608 2839 12610
rect 0 12552 2778 12608
rect 2834 12552 2839 12608
rect 0 12550 2839 12552
rect 0 12520 800 12550
rect 2773 12547 2839 12550
rect 15469 12610 15535 12613
rect 16062 12610 16068 12612
rect 15469 12608 16068 12610
rect 15469 12552 15474 12608
rect 15530 12552 16068 12608
rect 15469 12550 16068 12552
rect 15469 12547 15535 12550
rect 16062 12548 16068 12550
rect 16132 12548 16138 12612
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 10133 12474 10199 12477
rect 10501 12474 10567 12477
rect 16205 12476 16271 12477
rect 16205 12474 16252 12476
rect 10133 12472 10567 12474
rect 10133 12416 10138 12472
rect 10194 12416 10506 12472
rect 10562 12416 10567 12472
rect 10133 12414 10567 12416
rect 16160 12472 16252 12474
rect 16160 12416 16210 12472
rect 16160 12414 16252 12416
rect 10133 12411 10199 12414
rect 10501 12411 10567 12414
rect 16205 12412 16252 12414
rect 16316 12412 16322 12476
rect 17772 12474 17832 12686
rect 19200 12474 20000 12504
rect 17772 12414 20000 12474
rect 16205 12411 16271 12412
rect 19200 12384 20000 12414
rect 5257 12338 5323 12341
rect 9121 12338 9187 12341
rect 5257 12336 9187 12338
rect 5257 12280 5262 12336
rect 5318 12280 9126 12336
rect 9182 12280 9187 12336
rect 5257 12278 9187 12280
rect 5257 12275 5323 12278
rect 9121 12275 9187 12278
rect 10041 12338 10107 12341
rect 10358 12338 10364 12340
rect 10041 12336 10364 12338
rect 10041 12280 10046 12336
rect 10102 12280 10364 12336
rect 10041 12278 10364 12280
rect 10041 12275 10107 12278
rect 10358 12276 10364 12278
rect 10428 12276 10434 12340
rect 0 12202 800 12232
rect 4337 12202 4403 12205
rect 4981 12204 5047 12205
rect 4981 12202 5028 12204
rect 0 12200 4403 12202
rect 0 12144 4342 12200
rect 4398 12144 4403 12200
rect 0 12142 4403 12144
rect 4936 12200 5028 12202
rect 4936 12144 4986 12200
rect 4936 12142 5028 12144
rect 0 12112 800 12142
rect 4337 12139 4403 12142
rect 4981 12140 5028 12142
rect 5092 12140 5098 12204
rect 9622 12140 9628 12204
rect 9692 12202 9698 12204
rect 10225 12202 10291 12205
rect 9692 12200 10291 12202
rect 9692 12144 10230 12200
rect 10286 12144 10291 12200
rect 9692 12142 10291 12144
rect 9692 12140 9698 12142
rect 4981 12139 5047 12140
rect 10225 12139 10291 12142
rect 19200 12066 20000 12096
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 19152 11976 20000 12066
rect 3601 11930 3667 11933
rect 3601 11928 5274 11930
rect 3601 11872 3606 11928
rect 3662 11872 5274 11928
rect 3601 11870 5274 11872
rect 3601 11867 3667 11870
rect 0 11794 800 11824
rect 5073 11794 5139 11797
rect 0 11792 5139 11794
rect 0 11736 5078 11792
rect 5134 11736 5139 11792
rect 0 11734 5139 11736
rect 5214 11794 5274 11870
rect 19152 11828 19212 11976
rect 11145 11794 11211 11797
rect 5214 11792 11211 11794
rect 5214 11736 11150 11792
rect 11206 11736 11211 11792
rect 5214 11734 11211 11736
rect 0 11704 800 11734
rect 5073 11731 5139 11734
rect 11145 11731 11211 11734
rect 11462 11732 11468 11796
rect 11532 11794 11538 11796
rect 11697 11794 11763 11797
rect 13721 11796 13787 11797
rect 17953 11796 18019 11797
rect 11532 11792 11763 11794
rect 11532 11736 11702 11792
rect 11758 11736 11763 11792
rect 11532 11734 11763 11736
rect 11532 11732 11538 11734
rect 11697 11731 11763 11734
rect 13670 11732 13676 11796
rect 13740 11794 13787 11796
rect 13740 11792 13832 11794
rect 13782 11736 13832 11792
rect 13740 11734 13832 11736
rect 13740 11732 13787 11734
rect 17902 11732 17908 11796
rect 17972 11794 18019 11796
rect 18505 11794 18571 11797
rect 19060 11794 19212 11828
rect 17972 11792 18064 11794
rect 18014 11736 18064 11792
rect 17972 11734 18064 11736
rect 18505 11792 19212 11794
rect 18505 11736 18510 11792
rect 18566 11768 19212 11792
rect 18566 11736 19120 11768
rect 18505 11734 19120 11736
rect 17972 11732 18019 11734
rect 13721 11731 13787 11732
rect 17953 11731 18019 11732
rect 18505 11731 18571 11734
rect 1117 11658 1183 11661
rect 5349 11658 5415 11661
rect 1117 11656 5415 11658
rect 1117 11600 1122 11656
rect 1178 11600 5354 11656
rect 5410 11600 5415 11656
rect 1117 11598 5415 11600
rect 1117 11595 1183 11598
rect 5349 11595 5415 11598
rect 17493 11658 17559 11661
rect 19200 11658 20000 11688
rect 17493 11656 20000 11658
rect 17493 11600 17498 11656
rect 17554 11600 20000 11656
rect 17493 11598 20000 11600
rect 17493 11595 17559 11598
rect 19200 11568 20000 11598
rect 4429 11522 4495 11525
rect 7005 11522 7071 11525
rect 4429 11520 7071 11522
rect 4429 11464 4434 11520
rect 4490 11464 7010 11520
rect 7066 11464 7071 11520
rect 4429 11462 7071 11464
rect 4429 11459 4495 11462
rect 7005 11459 7071 11462
rect 3165 11456 3481 11457
rect 0 11386 800 11416
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 2865 11386 2931 11389
rect 0 11384 2931 11386
rect 0 11328 2870 11384
rect 2926 11328 2931 11384
rect 0 11326 2931 11328
rect 0 11296 800 11326
rect 2865 11323 2931 11326
rect 14457 11386 14523 11389
rect 14774 11386 14780 11388
rect 14457 11384 14780 11386
rect 14457 11328 14462 11384
rect 14518 11328 14780 11384
rect 14457 11326 14780 11328
rect 14457 11323 14523 11326
rect 14774 11324 14780 11326
rect 14844 11324 14850 11388
rect 4286 11188 4292 11252
rect 4356 11250 4362 11252
rect 11053 11250 11119 11253
rect 4356 11248 11119 11250
rect 4356 11192 11058 11248
rect 11114 11192 11119 11248
rect 4356 11190 11119 11192
rect 4356 11188 4362 11190
rect 11053 11187 11119 11190
rect 18321 11250 18387 11253
rect 19200 11250 20000 11280
rect 18321 11248 20000 11250
rect 18321 11192 18326 11248
rect 18382 11192 20000 11248
rect 18321 11190 20000 11192
rect 18321 11187 18387 11190
rect 19200 11160 20000 11190
rect 2037 11114 2103 11117
rect 7189 11114 7255 11117
rect 2037 11112 7255 11114
rect 2037 11056 2042 11112
rect 2098 11056 7194 11112
rect 7250 11056 7255 11112
rect 2037 11054 7255 11056
rect 2037 11051 2103 11054
rect 7189 11051 7255 11054
rect 0 10978 800 11008
rect 5165 10978 5231 10981
rect 0 10976 5231 10978
rect 0 10920 5170 10976
rect 5226 10920 5231 10976
rect 0 10918 5231 10920
rect 0 10888 800 10918
rect 5165 10915 5231 10918
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 19200 10842 20000 10872
rect 19152 10752 20000 10842
rect 2221 10706 2287 10709
rect 2497 10706 2563 10709
rect 2221 10704 2563 10706
rect 2221 10648 2226 10704
rect 2282 10648 2502 10704
rect 2558 10648 2563 10704
rect 2221 10646 2563 10648
rect 2221 10643 2287 10646
rect 2497 10643 2563 10646
rect 4429 10706 4495 10709
rect 5533 10706 5599 10709
rect 4429 10704 5599 10706
rect 4429 10648 4434 10704
rect 4490 10648 5538 10704
rect 5594 10648 5599 10704
rect 4429 10646 5599 10648
rect 4429 10643 4495 10646
rect 5533 10643 5599 10646
rect 8150 10644 8156 10708
rect 8220 10706 8226 10708
rect 8661 10706 8727 10709
rect 8220 10704 8727 10706
rect 8220 10648 8666 10704
rect 8722 10648 8727 10704
rect 8220 10646 8727 10648
rect 8220 10644 8226 10646
rect 8661 10643 8727 10646
rect 17677 10706 17743 10709
rect 19152 10706 19212 10752
rect 17677 10704 19212 10706
rect 17677 10648 17682 10704
rect 17738 10648 19212 10704
rect 17677 10646 19212 10648
rect 17677 10643 17743 10646
rect 0 10570 800 10600
rect 3969 10570 4035 10573
rect 0 10568 4035 10570
rect 0 10512 3974 10568
rect 4030 10512 4035 10568
rect 0 10510 4035 10512
rect 0 10480 800 10510
rect 3969 10507 4035 10510
rect 4521 10434 4587 10437
rect 5165 10434 5231 10437
rect 4521 10432 5231 10434
rect 4521 10376 4526 10432
rect 4582 10376 5170 10432
rect 5226 10376 5231 10432
rect 4521 10374 5231 10376
rect 4521 10371 4587 10374
rect 5165 10371 5231 10374
rect 18321 10434 18387 10437
rect 19200 10434 20000 10464
rect 18321 10432 20000 10434
rect 18321 10376 18326 10432
rect 18382 10376 20000 10432
rect 18321 10374 20000 10376
rect 18321 10371 18387 10374
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 19200 10344 20000 10374
rect 16482 10303 16798 10304
rect 9121 10300 9187 10301
rect 9070 10236 9076 10300
rect 9140 10298 9187 10300
rect 9140 10296 9232 10298
rect 9182 10240 9232 10296
rect 9140 10238 9232 10240
rect 9140 10236 9187 10238
rect 9121 10235 9187 10236
rect 0 10162 800 10192
rect 0 10102 2790 10162
rect 0 10072 800 10102
rect 2730 10026 2790 10102
rect 2957 10026 3023 10029
rect 2730 10024 3023 10026
rect 2730 9968 2962 10024
rect 3018 9968 3023 10024
rect 2730 9966 3023 9968
rect 2957 9963 3023 9966
rect 3877 10026 3943 10029
rect 4153 10026 4219 10029
rect 5441 10026 5507 10029
rect 3877 10024 4219 10026
rect 3877 9968 3882 10024
rect 3938 9968 4158 10024
rect 4214 9968 4219 10024
rect 3877 9966 4219 9968
rect 3877 9963 3943 9966
rect 4153 9963 4219 9966
rect 5260 10024 5507 10026
rect 5260 9968 5446 10024
rect 5502 9968 5507 10024
rect 5260 9966 5507 9968
rect 2497 9890 2563 9893
rect 5022 9890 5028 9892
rect 2497 9888 5028 9890
rect 2497 9832 2502 9888
rect 2558 9832 5028 9888
rect 2497 9830 5028 9832
rect 2497 9827 2563 9830
rect 5022 9828 5028 9830
rect 5092 9890 5098 9892
rect 5260 9890 5320 9966
rect 5441 9963 5507 9966
rect 18321 10026 18387 10029
rect 19200 10026 20000 10056
rect 18321 10024 20000 10026
rect 18321 9968 18326 10024
rect 18382 9968 20000 10024
rect 18321 9966 20000 9968
rect 18321 9963 18387 9966
rect 19200 9936 20000 9966
rect 5092 9830 5320 9890
rect 5092 9828 5098 9830
rect 5384 9824 5700 9825
rect 0 9754 800 9784
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 0 9694 5090 9754
rect 0 9664 800 9694
rect 4061 9618 4127 9621
rect 1350 9616 4127 9618
rect 1350 9560 4066 9616
rect 4122 9560 4127 9616
rect 1350 9558 4127 9560
rect 5030 9618 5090 9694
rect 5625 9618 5691 9621
rect 5030 9616 5691 9618
rect 5030 9560 5630 9616
rect 5686 9560 5691 9616
rect 5030 9558 5691 9560
rect 0 9346 800 9376
rect 1350 9346 1410 9558
rect 4061 9555 4127 9558
rect 5625 9555 5691 9558
rect 7046 9556 7052 9620
rect 7116 9618 7122 9620
rect 8661 9618 8727 9621
rect 7116 9616 8727 9618
rect 7116 9560 8666 9616
rect 8722 9560 8727 9616
rect 7116 9558 8727 9560
rect 7116 9556 7122 9558
rect 8661 9555 8727 9558
rect 9121 9618 9187 9621
rect 9254 9618 9260 9620
rect 9121 9616 9260 9618
rect 9121 9560 9126 9616
rect 9182 9560 9260 9616
rect 9121 9558 9260 9560
rect 9121 9555 9187 9558
rect 9254 9556 9260 9558
rect 9324 9556 9330 9620
rect 19200 9528 20000 9648
rect 2313 9482 2379 9485
rect 2865 9482 2931 9485
rect 2313 9480 2931 9482
rect 2313 9424 2318 9480
rect 2374 9424 2870 9480
rect 2926 9424 2931 9480
rect 2313 9422 2931 9424
rect 2313 9419 2379 9422
rect 2865 9419 2931 9422
rect 3417 9482 3483 9485
rect 4245 9482 4311 9485
rect 6637 9482 6703 9485
rect 3417 9480 6703 9482
rect 3417 9424 3422 9480
rect 3478 9424 4250 9480
rect 4306 9424 6642 9480
rect 6698 9424 6703 9480
rect 3417 9422 6703 9424
rect 3417 9419 3483 9422
rect 4245 9419 4311 9422
rect 6637 9419 6703 9422
rect 7414 9420 7420 9484
rect 7484 9482 7490 9484
rect 8109 9482 8175 9485
rect 7484 9480 8175 9482
rect 7484 9424 8114 9480
rect 8170 9424 8175 9480
rect 7484 9422 8175 9424
rect 7484 9420 7490 9422
rect 8109 9419 8175 9422
rect 0 9286 1410 9346
rect 4153 9346 4219 9349
rect 5257 9346 5323 9349
rect 4153 9344 5323 9346
rect 4153 9288 4158 9344
rect 4214 9288 5262 9344
rect 5318 9288 5323 9344
rect 4153 9286 5323 9288
rect 0 9256 800 9286
rect 4153 9283 4219 9286
rect 5257 9283 5323 9286
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 3693 9210 3759 9213
rect 4337 9210 4403 9213
rect 3693 9208 4403 9210
rect 3693 9152 3698 9208
rect 3754 9152 4342 9208
rect 4398 9152 4403 9208
rect 3693 9150 4403 9152
rect 3693 9147 3759 9150
rect 4337 9147 4403 9150
rect 5206 9148 5212 9212
rect 5276 9210 5282 9212
rect 5533 9210 5599 9213
rect 5276 9208 5599 9210
rect 5276 9152 5538 9208
rect 5594 9152 5599 9208
rect 5276 9150 5599 9152
rect 5276 9148 5282 9150
rect 5533 9147 5599 9150
rect 6678 9148 6684 9212
rect 6748 9210 6754 9212
rect 6821 9210 6887 9213
rect 6748 9208 6887 9210
rect 6748 9152 6826 9208
rect 6882 9152 6887 9208
rect 6748 9150 6887 9152
rect 6748 9148 6754 9150
rect 6821 9147 6887 9150
rect 18321 9210 18387 9213
rect 19200 9210 20000 9240
rect 18321 9208 20000 9210
rect 18321 9152 18326 9208
rect 18382 9152 20000 9208
rect 18321 9150 20000 9152
rect 18321 9147 18387 9150
rect 19200 9120 20000 9150
rect 2998 9012 3004 9076
rect 3068 9074 3074 9076
rect 6177 9074 6243 9077
rect 3068 9072 6243 9074
rect 3068 9016 6182 9072
rect 6238 9016 6243 9072
rect 3068 9014 6243 9016
rect 3068 9012 3074 9014
rect 6177 9011 6243 9014
rect 0 8938 800 8968
rect 3509 8938 3575 8941
rect 0 8936 3575 8938
rect 0 8880 3514 8936
rect 3570 8880 3575 8936
rect 0 8878 3575 8880
rect 0 8848 800 8878
rect 3509 8875 3575 8878
rect 19200 8805 20000 8832
rect 4245 8802 4311 8805
rect 4470 8802 4476 8804
rect 4245 8800 4476 8802
rect 4245 8744 4250 8800
rect 4306 8744 4476 8800
rect 4245 8742 4476 8744
rect 4245 8739 4311 8742
rect 4470 8740 4476 8742
rect 4540 8740 4546 8804
rect 19149 8800 20000 8805
rect 19149 8744 19154 8800
rect 19210 8744 20000 8800
rect 19149 8739 20000 8744
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 19200 8712 20000 8739
rect 18701 8671 19017 8672
rect 0 8530 800 8560
rect 4061 8530 4127 8533
rect 7189 8532 7255 8533
rect 7189 8530 7236 8532
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 7144 8528 7236 8530
rect 7144 8472 7194 8528
rect 7144 8470 7236 8472
rect 0 8440 800 8470
rect 4061 8467 4127 8470
rect 7189 8468 7236 8470
rect 7300 8468 7306 8532
rect 7189 8467 7255 8468
rect 19200 8304 20000 8424
rect 3165 8192 3481 8193
rect 0 8122 800 8152
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 2957 8122 3023 8125
rect 0 8120 3023 8122
rect 0 8064 2962 8120
rect 3018 8064 3023 8120
rect 0 8062 3023 8064
rect 0 8032 800 8062
rect 2957 8059 3023 8062
rect 4102 8060 4108 8124
rect 4172 8122 4178 8124
rect 5257 8122 5323 8125
rect 4172 8120 5323 8122
rect 4172 8064 5262 8120
rect 5318 8064 5323 8120
rect 4172 8062 5323 8064
rect 4172 8060 4178 8062
rect 5257 8059 5323 8062
rect 18321 7986 18387 7989
rect 19200 7986 20000 8016
rect 18321 7984 20000 7986
rect 18321 7928 18326 7984
rect 18382 7928 20000 7984
rect 18321 7926 20000 7928
rect 18321 7923 18387 7926
rect 19200 7896 20000 7926
rect 0 7714 800 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 800 7654
rect 4061 7651 4127 7654
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 19200 7578 20000 7608
rect 19152 7488 20000 7578
rect 5809 7442 5875 7445
rect 6126 7442 6132 7444
rect 5809 7440 6132 7442
rect 5809 7384 5814 7440
rect 5870 7384 6132 7440
rect 5809 7382 6132 7384
rect 5809 7379 5875 7382
rect 6126 7380 6132 7382
rect 6196 7380 6202 7444
rect 18321 7442 18387 7445
rect 19152 7442 19212 7488
rect 18321 7440 19212 7442
rect 18321 7384 18326 7440
rect 18382 7384 19212 7440
rect 18321 7382 19212 7384
rect 18321 7379 18387 7382
rect 0 7306 800 7336
rect 3969 7306 4035 7309
rect 0 7304 4035 7306
rect 0 7248 3974 7304
rect 4030 7248 4035 7304
rect 0 7246 4035 7248
rect 0 7216 800 7246
rect 3969 7243 4035 7246
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 19200 7080 20000 7200
rect 16482 7039 16798 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 18321 6762 18387 6765
rect 19200 6762 20000 6792
rect 18321 6760 20000 6762
rect 18321 6704 18326 6760
rect 18382 6704 20000 6760
rect 18321 6702 20000 6704
rect 18321 6699 18387 6702
rect 19200 6672 20000 6702
rect 5384 6560 5700 6561
rect 0 6490 800 6520
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 2865 6490 2931 6493
rect 0 6488 2931 6490
rect 0 6432 2870 6488
rect 2926 6432 2931 6488
rect 0 6430 2931 6432
rect 0 6400 800 6430
rect 2865 6427 2931 6430
rect 18321 6354 18387 6357
rect 19200 6354 20000 6384
rect 18321 6352 20000 6354
rect 18321 6296 18326 6352
rect 18382 6296 20000 6352
rect 18321 6294 20000 6296
rect 18321 6291 18387 6294
rect 19200 6264 20000 6294
rect 0 6082 800 6112
rect 2957 6082 3023 6085
rect 0 6080 3023 6082
rect 0 6024 2962 6080
rect 3018 6024 3023 6080
rect 0 6022 3023 6024
rect 0 5992 800 6022
rect 2957 6019 3023 6022
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 19200 5856 20000 5976
rect 0 5674 800 5704
rect 3969 5674 4035 5677
rect 0 5672 4035 5674
rect 0 5616 3974 5672
rect 4030 5616 4035 5672
rect 0 5614 4035 5616
rect 0 5584 800 5614
rect 3969 5611 4035 5614
rect 18321 5674 18387 5677
rect 18321 5672 19212 5674
rect 18321 5616 18326 5672
rect 18382 5616 19212 5672
rect 18321 5614 19212 5616
rect 18321 5611 18387 5614
rect 19152 5568 19212 5614
rect 19152 5478 20000 5568
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 19200 5448 20000 5478
rect 18701 5407 19017 5408
rect 0 5266 800 5296
rect 1577 5266 1643 5269
rect 0 5264 1643 5266
rect 0 5208 1582 5264
rect 1638 5208 1643 5264
rect 0 5206 1643 5208
rect 0 5176 800 5206
rect 1577 5203 1643 5206
rect 18321 5130 18387 5133
rect 19200 5130 20000 5160
rect 18321 5128 20000 5130
rect 18321 5072 18326 5128
rect 18382 5072 20000 5128
rect 18321 5070 20000 5072
rect 18321 5067 18387 5070
rect 19200 5040 20000 5070
rect 3165 4928 3481 4929
rect 0 4768 800 4888
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 19200 4632 20000 4752
rect 0 4450 800 4480
rect 1669 4450 1735 4453
rect 0 4448 1735 4450
rect 0 4392 1674 4448
rect 1730 4392 1735 4448
rect 0 4390 1735 4392
rect 0 4360 800 4390
rect 1669 4387 1735 4390
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 19200 4317 20000 4344
rect 19149 4312 20000 4317
rect 19149 4256 19154 4312
rect 19210 4256 20000 4312
rect 19149 4251 20000 4256
rect 19200 4224 20000 4251
rect 0 4042 800 4072
rect 1577 4042 1643 4045
rect 0 4040 1643 4042
rect 0 3984 1582 4040
rect 1638 3984 1643 4040
rect 0 3982 1643 3984
rect 0 3952 800 3982
rect 1577 3979 1643 3982
rect 18321 3906 18387 3909
rect 19200 3906 20000 3936
rect 18321 3904 20000 3906
rect 18321 3848 18326 3904
rect 18382 3848 20000 3904
rect 18321 3846 20000 3848
rect 18321 3843 18387 3846
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 19200 3816 20000 3846
rect 16482 3775 16798 3776
rect 0 3544 800 3664
rect 19200 3408 20000 3528
rect 5384 3296 5700 3297
rect 0 3226 800 3256
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 1577 3226 1643 3229
rect 0 3224 1643 3226
rect 0 3168 1582 3224
rect 1638 3168 1643 3224
rect 0 3166 1643 3168
rect 0 3136 800 3166
rect 1577 3163 1643 3166
rect 18321 3090 18387 3093
rect 19200 3090 20000 3120
rect 18321 3088 20000 3090
rect 18321 3032 18326 3088
rect 18382 3032 20000 3088
rect 18321 3030 20000 3032
rect 18321 3027 18387 3030
rect 19200 3000 20000 3030
rect 0 2818 800 2848
rect 1577 2818 1643 2821
rect 0 2816 1643 2818
rect 0 2760 1582 2816
rect 1638 2760 1643 2816
rect 0 2758 1643 2760
rect 0 2728 800 2758
rect 1577 2755 1643 2758
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 18321 2682 18387 2685
rect 19200 2682 20000 2712
rect 18321 2680 20000 2682
rect 18321 2624 18326 2680
rect 18382 2624 20000 2680
rect 18321 2622 20000 2624
rect 18321 2619 18387 2622
rect 19200 2592 20000 2622
rect 0 2320 800 2440
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 19200 2184 20000 2304
rect 18701 2143 19017 2144
rect 0 2002 800 2032
rect 2221 2002 2287 2005
rect 0 2000 2287 2002
rect 0 1944 2226 2000
rect 2282 1944 2287 2000
rect 0 1942 2287 1944
rect 0 1912 800 1942
rect 2221 1939 2287 1942
rect 18321 1866 18387 1869
rect 19200 1866 20000 1896
rect 18321 1864 20000 1866
rect 18321 1808 18326 1864
rect 18382 1808 20000 1864
rect 18321 1806 20000 1808
rect 18321 1803 18387 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
rect 17677 1458 17743 1461
rect 19200 1458 20000 1488
rect 17677 1456 20000 1458
rect 17677 1400 17682 1456
rect 17738 1400 20000 1456
rect 17677 1398 20000 1400
rect 17677 1395 17743 1398
rect 19200 1368 20000 1398
rect 19200 960 20000 1080
<< via3 >>
rect 7236 18532 7300 18596
rect 13676 18532 13740 18596
rect 6132 18260 6196 18324
rect 9260 17852 9324 17916
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 7420 17172 7484 17236
rect 14780 17172 14844 17236
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 11468 17036 11532 17100
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 10364 16628 10428 16692
rect 9076 16492 9140 16556
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 4292 16220 4356 16284
rect 8156 16084 8220 16148
rect 5212 15948 5276 16012
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 7052 15540 7116 15604
rect 9628 15540 9692 15604
rect 10548 15404 10612 15468
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 15884 14996 15948 15060
rect 16252 14996 16316 15060
rect 4476 14724 4540 14788
rect 16068 14724 16132 14788
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 3004 14588 3068 14652
rect 17908 14316 17972 14380
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 4108 13908 4172 13972
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 6684 13500 6748 13564
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 10548 12820 10612 12884
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 15884 13092 15948 13156
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 16068 12548 16132 12612
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 16252 12472 16316 12476
rect 16252 12416 16266 12472
rect 16266 12416 16316 12472
rect 16252 12412 16316 12416
rect 10364 12276 10428 12340
rect 5028 12200 5092 12204
rect 5028 12144 5042 12200
rect 5042 12144 5092 12200
rect 5028 12140 5092 12144
rect 9628 12140 9692 12204
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 11468 11732 11532 11796
rect 13676 11792 13740 11796
rect 13676 11736 13726 11792
rect 13726 11736 13740 11792
rect 13676 11732 13740 11736
rect 17908 11792 17972 11796
rect 17908 11736 17958 11792
rect 17958 11736 17972 11792
rect 17908 11732 17972 11736
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 14780 11324 14844 11388
rect 4292 11188 4356 11252
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 8156 10644 8220 10708
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 9076 10296 9140 10300
rect 9076 10240 9126 10296
rect 9126 10240 9140 10296
rect 9076 10236 9140 10240
rect 5028 9828 5092 9892
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 7052 9556 7116 9620
rect 9260 9556 9324 9620
rect 7420 9420 7484 9484
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5212 9148 5276 9212
rect 6684 9148 6748 9212
rect 3004 9012 3068 9076
rect 4476 8740 4540 8804
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 7236 8528 7300 8532
rect 7236 8472 7250 8528
rect 7250 8472 7300 8528
rect 7236 8468 7300 8472
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 4108 8060 4172 8124
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 6132 7380 6196 7444
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 7235 18596 7301 18597
rect 7235 18532 7236 18596
rect 7300 18532 7301 18596
rect 7235 18531 7301 18532
rect 13675 18596 13741 18597
rect 13675 18532 13676 18596
rect 13740 18532 13741 18596
rect 13675 18531 13741 18532
rect 6131 18324 6197 18325
rect 6131 18260 6132 18324
rect 6196 18260 6197 18324
rect 6131 18259 6197 18260
rect 3163 16896 3483 17456
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 5382 17440 5702 17456
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 4291 16284 4357 16285
rect 4291 16220 4292 16284
rect 4356 16220 4357 16284
rect 4291 16219 4357 16220
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3003 14652 3069 14653
rect 3003 14588 3004 14652
rect 3068 14588 3069 14652
rect 3003 14587 3069 14588
rect 3006 9077 3066 14587
rect 3163 13632 3483 14656
rect 4107 13972 4173 13973
rect 4107 13908 4108 13972
rect 4172 13908 4173 13972
rect 4107 13907 4173 13908
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3003 9076 3069 9077
rect 3003 9012 3004 9076
rect 3068 9012 3069 9076
rect 3003 9011 3069 9012
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 4110 8125 4170 13907
rect 4294 11253 4354 16219
rect 5211 16012 5277 16013
rect 5211 15948 5212 16012
rect 5276 15948 5277 16012
rect 5211 15947 5277 15948
rect 4475 14788 4541 14789
rect 4475 14724 4476 14788
rect 4540 14724 4541 14788
rect 4475 14723 4541 14724
rect 4291 11252 4357 11253
rect 4291 11188 4292 11252
rect 4356 11188 4357 11252
rect 4291 11187 4357 11188
rect 4478 8805 4538 14723
rect 5027 12204 5093 12205
rect 5027 12140 5028 12204
rect 5092 12140 5093 12204
rect 5027 12139 5093 12140
rect 5030 9893 5090 12139
rect 5027 9892 5093 9893
rect 5027 9828 5028 9892
rect 5092 9828 5093 9892
rect 5027 9827 5093 9828
rect 5214 9213 5274 15947
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5211 9212 5277 9213
rect 5211 9148 5212 9212
rect 5276 9148 5277 9212
rect 5211 9147 5277 9148
rect 4475 8804 4541 8805
rect 4475 8740 4476 8804
rect 4540 8740 4541 8804
rect 4475 8739 4541 8740
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 4107 8124 4173 8125
rect 4107 8060 4108 8124
rect 4172 8060 4173 8124
rect 4107 8059 4173 8060
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 6134 7445 6194 18259
rect 7051 15604 7117 15605
rect 7051 15540 7052 15604
rect 7116 15540 7117 15604
rect 7051 15539 7117 15540
rect 6683 13564 6749 13565
rect 6683 13500 6684 13564
rect 6748 13500 6749 13564
rect 6683 13499 6749 13500
rect 6686 9213 6746 13499
rect 7054 9621 7114 15539
rect 7051 9620 7117 9621
rect 7051 9556 7052 9620
rect 7116 9556 7117 9620
rect 7051 9555 7117 9556
rect 6683 9212 6749 9213
rect 6683 9148 6684 9212
rect 6748 9148 6749 9212
rect 6683 9147 6749 9148
rect 7238 8533 7298 18531
rect 9259 17916 9325 17917
rect 9259 17852 9260 17916
rect 9324 17852 9325 17916
rect 9259 17851 9325 17852
rect 7419 17236 7485 17237
rect 7419 17172 7420 17236
rect 7484 17172 7485 17236
rect 7419 17171 7485 17172
rect 7422 9485 7482 17171
rect 7602 16896 7922 17456
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 9075 16556 9141 16557
rect 9075 16492 9076 16556
rect 9140 16492 9141 16556
rect 9075 16491 9141 16492
rect 8155 16148 8221 16149
rect 8155 16084 8156 16148
rect 8220 16084 8221 16148
rect 8155 16083 8221 16084
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 8158 10709 8218 16083
rect 8155 10708 8221 10709
rect 8155 10644 8156 10708
rect 8220 10644 8221 10708
rect 8155 10643 8221 10644
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7419 9484 7485 9485
rect 7419 9420 7420 9484
rect 7484 9420 7485 9484
rect 7419 9419 7485 9420
rect 7602 9280 7922 10304
rect 9078 10301 9138 16491
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 9262 9621 9322 17851
rect 9821 17440 10141 17456
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 11467 17100 11533 17101
rect 11467 17036 11468 17100
rect 11532 17036 11533 17100
rect 11467 17035 11533 17036
rect 10363 16692 10429 16693
rect 10363 16628 10364 16692
rect 10428 16628 10429 16692
rect 10363 16627 10429 16628
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9627 15604 9693 15605
rect 9627 15540 9628 15604
rect 9692 15540 9693 15604
rect 9627 15539 9693 15540
rect 9630 12205 9690 15539
rect 9821 15264 10141 16288
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9627 12204 9693 12205
rect 9627 12140 9628 12204
rect 9692 12140 9693 12204
rect 9627 12139 9693 12140
rect 9821 12000 10141 13024
rect 10366 12341 10426 16627
rect 10547 15468 10613 15469
rect 10547 15404 10548 15468
rect 10612 15404 10613 15468
rect 10547 15403 10613 15404
rect 10550 12885 10610 15403
rect 10547 12884 10613 12885
rect 10547 12820 10548 12884
rect 10612 12820 10613 12884
rect 10547 12819 10613 12820
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 11470 11797 11530 17035
rect 12041 16896 12361 17456
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 14720 12361 15744
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 11467 11796 11533 11797
rect 11467 11732 11468 11796
rect 11532 11732 11533 11796
rect 11467 11731 11533 11732
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9259 9620 9325 9621
rect 9259 9556 9260 9620
rect 9324 9556 9325 9620
rect 9259 9555 9325 9556
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7235 8532 7301 8533
rect 7235 8468 7236 8532
rect 7300 8468 7301 8532
rect 7235 8467 7301 8468
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 6131 7444 6197 7445
rect 6131 7380 6132 7444
rect 6196 7380 6197 7444
rect 6131 7379 6197 7380
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 11456 12361 12480
rect 13678 11797 13738 18531
rect 14260 17440 14580 17456
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14779 17236 14845 17237
rect 14779 17172 14780 17236
rect 14844 17172 14845 17236
rect 14779 17171 14845 17172
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 14260 15264 14580 16288
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 10912 14580 11936
rect 14782 11389 14842 17171
rect 16480 16896 16800 17456
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 15883 15060 15949 15061
rect 15883 14996 15884 15060
rect 15948 14996 15949 15060
rect 15883 14995 15949 14996
rect 16251 15060 16317 15061
rect 16251 14996 16252 15060
rect 16316 14996 16317 15060
rect 16251 14995 16317 14996
rect 15886 13157 15946 14995
rect 16067 14788 16133 14789
rect 16067 14724 16068 14788
rect 16132 14724 16133 14788
rect 16067 14723 16133 14724
rect 15883 13156 15949 13157
rect 15883 13092 15884 13156
rect 15948 13092 15949 13156
rect 15883 13091 15949 13092
rect 16070 12613 16130 14723
rect 16067 12612 16133 12613
rect 16067 12548 16068 12612
rect 16132 12548 16133 12612
rect 16067 12547 16133 12548
rect 16254 12477 16314 14995
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 18699 17440 19019 17456
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 17907 14380 17973 14381
rect 17907 14316 17908 14380
rect 17972 14316 17973 14380
rect 17907 14315 17973 14316
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16251 12476 16317 12477
rect 16251 12412 16252 12476
rect 16316 12412 16317 12476
rect 16251 12411 16317 12412
rect 16480 11456 16800 12480
rect 17910 11797 17970 14315
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 17907 11796 17973 11797
rect 17907 11732 17908 11796
rect 17972 11732 17973 11796
rect 17907 11731 17973 11732
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 14779 11388 14845 11389
rect 14779 11324 14780 11388
rect 14844 11324 14845 11388
rect 14779 11323 14845 11324
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 16192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1666464484
transform -1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1666464484
transform -1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1666464484
transform -1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1666464484
transform -1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1666464484
transform -1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1666464484
transform -1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1666464484
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1666464484
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1666464484
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1666464484
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1666464484
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1666464484
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_22
timestamp 1666464484
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_34
timestamp 1666464484
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1666464484
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1666464484
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1666464484
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1666464484
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1666464484
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1666464484
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_40
timestamp 1666464484
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_52
timestamp 1666464484
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_64
timestamp 1666464484
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1666464484
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp 1666464484
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp 1666464484
transform 1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_29
timestamp 1666464484
transform 1 0 3772 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1666464484
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1666464484
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1666464484
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1666464484
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1666464484
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1666464484
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1666464484
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1666464484
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_55
timestamp 1666464484
transform 1 0 6164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_67
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1666464484
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1666464484
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_10
timestamp 1666464484
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1666464484
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1666464484
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1666464484
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1666464484
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1666464484
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1666464484
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_61
timestamp 1666464484
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_67
timestamp 1666464484
transform 1 0 7268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_79
timestamp 1666464484
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1666464484
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1666464484
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1666464484
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1666464484
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1666464484
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1666464484
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1666464484
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1666464484
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1666464484
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_68
timestamp 1666464484
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1666464484
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1666464484
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1666464484
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1666464484
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1666464484
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1666464484
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1666464484
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1666464484
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_75
timestamp 1666464484
transform 1 0 8004 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_87
timestamp 1666464484
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_99
timestamp 1666464484
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1666464484
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1666464484
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1666464484
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1666464484
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1666464484
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1666464484
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1666464484
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1666464484
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_89
timestamp 1666464484
transform 1 0 9292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_101
timestamp 1666464484
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_113
timestamp 1666464484
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_125
timestamp 1666464484
transform 1 0 12604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1666464484
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1666464484
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1666464484
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1666464484
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_176
timestamp 1666464484
transform 1 0 17296 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_184
timestamp 1666464484
transform 1 0 18032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1666464484
transform 1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1666464484
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1666464484
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1666464484
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_76
timestamp 1666464484
transform 1 0 8096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1666464484
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_90
timestamp 1666464484
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_96
timestamp 1666464484
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1666464484
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1666464484
transform 1 0 15548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_160
timestamp 1666464484
transform 1 0 15824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1666464484
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1666464484
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_39
timestamp 1666464484
transform 1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_48
timestamp 1666464484
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1666464484
transform 1 0 6348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1666464484
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_71
timestamp 1666464484
transform 1 0 7636 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1666464484
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1666464484
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_96
timestamp 1666464484
transform 1 0 9936 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_108
timestamp 1666464484
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_120
timestamp 1666464484
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1666464484
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1666464484
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1666464484
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1666464484
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1666464484
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1666464484
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_26
timestamp 1666464484
transform 1 0 3496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1666464484
transform 1 0 5336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1666464484
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_64
timestamp 1666464484
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1666464484
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1666464484
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1666464484
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1666464484
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1666464484
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1666464484
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1666464484
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1666464484
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1666464484
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1666464484
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_38
timestamp 1666464484
transform 1 0 4600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1666464484
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1666464484
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1666464484
transform 1 0 6900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1666464484
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1666464484
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1666464484
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1666464484
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_117
timestamp 1666464484
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_129
timestamp 1666464484
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1666464484
transform 1 0 13524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1666464484
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1666464484
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1666464484
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1666464484
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1666464484
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1666464484
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1666464484
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1666464484
transform 1 0 4968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_61
timestamp 1666464484
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1666464484
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_72
timestamp 1666464484
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_76
timestamp 1666464484
transform 1 0 8096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1666464484
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1666464484
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1666464484
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1666464484
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1666464484
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_118
timestamp 1666464484
transform 1 0 11960 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_126
timestamp 1666464484
transform 1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1666464484
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_138
timestamp 1666464484
transform 1 0 13800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1666464484
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1666464484
transform 1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1666464484
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1666464484
transform 1 0 17572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1666464484
transform 1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_36
timestamp 1666464484
transform 1 0 4416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1666464484
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1666464484
transform 1 0 6072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1666464484
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1666464484
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1666464484
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1666464484
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1666464484
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1666464484
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1666464484
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_119
timestamp 1666464484
transform 1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1666464484
transform 1 0 12788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1666464484
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1666464484
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1666464484
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1666464484
transform 1 0 14812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1666464484
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1666464484
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1666464484
transform 1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1666464484
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1666464484
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1666464484
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_40
timestamp 1666464484
transform 1 0 4784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_46
timestamp 1666464484
transform 1 0 5336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1666464484
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_75
timestamp 1666464484
transform 1 0 8004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_83
timestamp 1666464484
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1666464484
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1666464484
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1666464484
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1666464484
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1666464484
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1666464484
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1666464484
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1666464484
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1666464484
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1666464484
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1666464484
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1666464484
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp 1666464484
transform 1 0 4416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1666464484
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_54
timestamp 1666464484
transform 1 0 6072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_63
timestamp 1666464484
transform 1 0 6900 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_69
timestamp 1666464484
transform 1 0 7452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1666464484
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1666464484
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1666464484
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_120
timestamp 1666464484
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1666464484
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1666464484
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1666464484
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1666464484
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1666464484
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1666464484
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1666464484
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_31
timestamp 1666464484
transform 1 0 3956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1666464484
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1666464484
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1666464484
transform 1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_79
timestamp 1666464484
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1666464484
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_122
timestamp 1666464484
transform 1 0 12328 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1666464484
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1666464484
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_141
timestamp 1666464484
transform 1 0 14076 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1666464484
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1666464484
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1666464484
transform 1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1666464484
transform 1 0 18400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1666464484
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_47
timestamp 1666464484
transform 1 0 5428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_56
timestamp 1666464484
transform 1 0 6256 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_60
timestamp 1666464484
transform 1 0 6624 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1666464484
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_95
timestamp 1666464484
transform 1 0 9844 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1666464484
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_126
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_146
timestamp 1666464484
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_155
timestamp 1666464484
transform 1 0 15364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1666464484
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1666464484
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1666464484
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1666464484
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1666464484
transform 1 0 5152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1666464484
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1666464484
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_67
timestamp 1666464484
transform 1 0 7268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1666464484
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_87
timestamp 1666464484
transform 1 0 9108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_102
timestamp 1666464484
transform 1 0 10488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_120
timestamp 1666464484
transform 1 0 12144 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1666464484
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1666464484
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1666464484
transform 1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1666464484
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1666464484
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1666464484
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_71
timestamp 1666464484
transform 1 0 7636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1666464484
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 1666464484
transform 1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_113
timestamp 1666464484
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1666464484
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1666464484
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1666464484
transform 1 0 14536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1666464484
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1666464484
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1666464484
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1666464484
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1666464484
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1666464484
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1666464484
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1666464484
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1666464484
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1666464484
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1666464484
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_131
timestamp 1666464484
transform 1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1666464484
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1666464484
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1666464484
transform 1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_48
timestamp 1666464484
transform 1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_54
timestamp 1666464484
transform 1 0 6072 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1666464484
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1666464484
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1666464484
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1666464484
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_21
timestamp 1666464484
transform 1 0 3036 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1666464484
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1666464484
transform 1 0 4508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_43
timestamp 1666464484
transform 1 0 5060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1666464484
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1666464484
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1666464484
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1666464484
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1666464484
transform 1 0 13156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1666464484
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1666464484
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1666464484
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1666464484
transform 1 0 18400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _153_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3772 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _155_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1666464484
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _157_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4968 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _158_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2576 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _159_
timestamp 1666464484
transform -1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _160_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _162_
timestamp 1666464484
transform -1 0 4048 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _163_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _164_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _165_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3496 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _166_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5428 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _167_
timestamp 1666464484
transform -1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _168_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _169_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4416 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _170_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _171_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1666464484
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1666464484
transform -1 0 3036 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 1666464484
transform 1 0 2576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _175_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1666464484
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _177_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3496 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _178_
timestamp 1666464484
transform 1 0 5060 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _179_
timestamp 1666464484
transform -1 0 4600 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1666464484
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1666464484
transform -1 0 5244 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _182_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _183_
timestamp 1666464484
transform 1 0 1564 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1666464484
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _185_
timestamp 1666464484
transform 1 0 5336 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _186_
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _187_
timestamp 1666464484
transform -1 0 5796 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _189_
timestamp 1666464484
transform 1 0 3496 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1666464484
transform -1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _191_
timestamp 1666464484
transform -1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1666464484
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _193_
timestamp 1666464484
transform 1 0 5612 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _194_
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _195_
timestamp 1666464484
transform 1 0 6440 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1666464484
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 1666464484
transform 1 0 5612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _198_
timestamp 1666464484
transform -1 0 3956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _199_
timestamp 1666464484
transform -1 0 4600 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1666464484
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 1666464484
transform -1 0 6256 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _202_
timestamp 1666464484
transform 1 0 4324 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _203_
timestamp 1666464484
transform 1 0 4416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1666464484
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 1666464484
transform 1 0 5520 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 1666464484
transform -1 0 5244 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _207_
timestamp 1666464484
transform 1 0 1564 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1666464484
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _209_
timestamp 1666464484
transform -1 0 5428 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1666464484
transform -1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1666464484
transform 1 0 4324 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1666464484
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _213_
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1666464484
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _215_
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1666464484
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _217_
timestamp 1666464484
transform -1 0 12328 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1666464484
transform 1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _219_
timestamp 1666464484
transform -1 0 8096 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1666464484
transform 1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _221_
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _223_
timestamp 1666464484
transform 1 0 6164 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1666464484
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _225_
timestamp 1666464484
transform -1 0 9292 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 1666464484
transform -1 0 7820 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _227_
timestamp 1666464484
transform 1 0 5428 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1666464484
transform 1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _229_
timestamp 1666464484
transform -1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _230_
timestamp 1666464484
transform 1 0 6808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _231_
timestamp 1666464484
transform 1 0 6716 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1666464484
transform -1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _233_
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _234_
timestamp 1666464484
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _235_
timestamp 1666464484
transform -1 0 12144 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1666464484
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1666464484
transform -1 0 13156 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1666464484
transform -1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_
timestamp 1666464484
transform -1 0 17388 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1666464484
transform -1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _241_
timestamp 1666464484
transform 1 0 14904 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1666464484
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _243_
timestamp 1666464484
transform -1 0 18308 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1666464484
transform 1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _245_
timestamp 1666464484
transform -1 0 14444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _246_
timestamp 1666464484
transform 1 0 17848 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _247_
timestamp 1666464484
transform 1 0 15916 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1666464484
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1666464484
transform 1 0 16100 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1666464484
transform -1 0 13616 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _251_
timestamp 1666464484
transform -1 0 17296 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1666464484
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _253_
timestamp 1666464484
transform 1 0 15088 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _254_
timestamp 1666464484
transform -1 0 15732 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _255_
timestamp 1666464484
transform -1 0 18400 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1666464484
transform -1 0 13156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _257_
timestamp 1666464484
transform -1 0 18400 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1666464484
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _259_
timestamp 1666464484
transform -1 0 17480 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform -1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _261_
timestamp 1666464484
transform -1 0 16376 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform -1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _263_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11500 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1666464484
transform -1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1666464484
transform -1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _267_
timestamp 1666464484
transform -1 0 15548 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _269_
timestamp 1666464484
transform 1 0 15732 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _270_
timestamp 1666464484
transform 1 0 17848 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _271_
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1666464484
transform -1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1666464484
transform -1 0 13156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _274_
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _275_
timestamp 1666464484
transform 1 0 13892 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _276_
timestamp 1666464484
transform -1 0 17480 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _277_
timestamp 1666464484
transform -1 0 18400 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _278_
timestamp 1666464484
transform -1 0 12328 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1666464484
transform -1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _281_
timestamp 1666464484
transform -1 0 8648 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1666464484
transform -1 0 6808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _283_
timestamp 1666464484
transform -1 0 11500 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1666464484
transform -1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _285_
timestamp 1666464484
transform -1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _286_
timestamp 1666464484
transform -1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1666464484
transform 1 0 13064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _288_
timestamp 1666464484
transform 1 0 10580 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _289_
timestamp 1666464484
transform 1 0 7728 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _290_
timestamp 1666464484
transform 1 0 9292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _291_
timestamp 1666464484
transform -1 0 11040 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _292_
timestamp 1666464484
transform -1 0 9108 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1666464484
transform 1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1666464484
transform 1 0 8004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _295_
timestamp 1666464484
transform 1 0 3404 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1666464484
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _297_
timestamp 1666464484
transform -1 0 4508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _298_
timestamp 1666464484
transform -1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _299_
timestamp 1666464484
transform -1 0 5980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _300_
timestamp 1666464484
transform -1 0 4140 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1666464484
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _302_
timestamp 1666464484
transform -1 0 5152 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _303_
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _304_
timestamp 1666464484
transform -1 0 6348 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _305_
timestamp 1666464484
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _306_
timestamp 1666464484
transform 1 0 5244 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _307_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12052 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp 1666464484
transform 1 0 8464 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp 1666464484
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _311_
timestamp 1666464484
transform 1 0 1564 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _312_
timestamp 1666464484
transform 1 0 1564 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _313_
timestamp 1666464484
transform 1 0 1564 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _314_
timestamp 1666464484
transform 1 0 1564 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _315_
timestamp 1666464484
transform -1 0 3036 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _316_
timestamp 1666464484
transform 1 0 1564 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _317_
timestamp 1666464484
transform -1 0 5336 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _318_
timestamp 1666464484
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _319_
timestamp 1666464484
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _320_
timestamp 1666464484
transform 1 0 3956 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _321_
timestamp 1666464484
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _322_
timestamp 1666464484
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _323_
timestamp 1666464484
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _324_
timestamp 1666464484
transform -1 0 3036 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _325_
timestamp 1666464484
transform 1 0 8740 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1666464484
transform 1 0 7176 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1666464484
transform -1 0 10580 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1666464484
transform -1 0 8648 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1666464484
transform 1 0 10948 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1666464484
transform -1 0 10580 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1666464484
transform 1 0 11684 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1666464484
transform 1 0 16928 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1666464484
transform -1 0 16100 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1666464484
transform 1 0 16928 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _335_
timestamp 1666464484
transform 1 0 14904 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _336_
timestamp 1666464484
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _337_
timestamp 1666464484
transform 1 0 16928 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _338_
timestamp 1666464484
transform 1 0 16928 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1666464484
transform 1 0 6072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout31
timestamp 1666464484
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1666464484
transform -1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform 1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform -1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1666464484
transform -1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1666464484
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1666464484
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1666464484
transform 1 0 8464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1666464484
transform -1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1666464484
transform -1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1666464484
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1666464484
transform 1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1666464484
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1666464484
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1666464484
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1666464484
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1666464484
transform 1 0 17480 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1666464484
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform 1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform 1 0 17296 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform 1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform 1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform 1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform -1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform -1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform -1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform -1 0 5520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform -1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform -1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform -1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform -1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform -1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform -1 0 6992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform -1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_78
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_79
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_80
timestamp 1666464484
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_81
timestamp 1666464484
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_82
timestamp 1666464484
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_83
timestamp 1666464484
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_84
timestamp 1666464484
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_85
timestamp 1666464484
transform 1 0 13524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_86
timestamp 1666464484
transform 1 0 12880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_87
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_88
timestamp 1666464484
transform -1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_89
timestamp 1666464484
transform -1 0 12788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_90
timestamp 1666464484
transform -1 0 13800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_91
timestamp 1666464484
transform -1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_92
timestamp 1666464484
transform -1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_93
timestamp 1666464484
transform -1 0 8924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_94
timestamp 1666464484
transform -1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_95
timestamp 1666464484
transform -1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_96
timestamp 1666464484
transform -1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_97
timestamp 1666464484
transform -1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_98
timestamp 1666464484
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_99
timestamp 1666464484
transform -1 0 12144 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_100
timestamp 1666464484
transform -1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_101
timestamp 1666464484
transform -1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_102
timestamp 1666464484
transform -1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_103
timestamp 1666464484
transform -1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_104
timestamp 1666464484
transform -1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_105
timestamp 1666464484
transform -1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_106
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_107
timestamp 1666464484
transform -1 0 2484 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 19200 16872 20000 16992 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 19200 18096 20000 18216 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 19522 19200 19578 20000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 17314 19200 17370 20000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 15106 19200 15162 20000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 12898 19200 12954 20000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 10690 19200 10746 20000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 8482 19200 8538 20000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 6274 19200 6330 20000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 4066 19200 4122 20000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 1858 19200 1914 20000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 19200 17688 20000 17808 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 19200 18912 20000 19032 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 18050 19200 18106 20000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 15842 19200 15898 20000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 13634 19200 13690 20000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 11426 19200 11482 20000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 9218 19200 9274 20000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 7010 19200 7066 20000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 4802 19200 4858 20000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 2594 19200 2650 20000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 386 19200 442 20000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 19200 17280 20000 17400 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 18786 19200 18842 20000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 16578 19200 16634 20000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 14370 19200 14426 20000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 12162 19200 12218 20000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 7746 19200 7802 20000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 5538 19200 5594 20000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 3330 19200 3386 20000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 1122 19200 1178 20000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 3163 2128 3483 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7602 2128 7922 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 12041 2128 12361 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 16480 2128 16800 17456 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 5382 2128 5702 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 17456 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 9982 16864 9982 16864 0 vccd1
rlabel via1 10061 17408 10061 17408 0 vssd1
rlabel metal2 11730 14178 11730 14178 0 _000_
rlabel metal1 8678 13974 8678 13974 0 _001_
rlabel metal1 6072 13770 6072 13770 0 _002_
rlabel metal1 6256 12682 6256 12682 0 _003_
rlabel metal2 2254 8296 2254 8296 0 _004_
rlabel metal1 2300 7514 2300 7514 0 _005_
rlabel metal1 4646 9350 4646 9350 0 _006_
rlabel metal1 1840 6630 1840 6630 0 _007_
rlabel metal1 2990 7514 2990 7514 0 _008_
rlabel metal2 1794 9248 1794 9248 0 _009_
rlabel metal2 5198 9333 5198 9333 0 _010_
rlabel metal1 1416 17170 1416 17170 0 _011_
rlabel metal2 11822 12546 11822 12546 0 _012_
rlabel metal1 1564 6154 1564 6154 0 _013_
rlabel metal1 2065 16082 2065 16082 0 _014_
rlabel metal1 2111 14994 2111 14994 0 _015_
rlabel metal1 2318 14314 2318 14314 0 _016_
rlabel metal2 3358 16320 3358 16320 0 _017_
rlabel via1 9057 16082 9057 16082 0 _018_
rlabel metal1 7590 13192 7590 13192 0 _019_
rlabel metal1 10304 12954 10304 12954 0 _020_
rlabel metal1 8694 17102 8694 17102 0 _021_
rlabel metal1 11357 16490 11357 16490 0 _022_
rlabel metal1 10948 12954 10948 12954 0 _023_
rlabel metal1 11536 17170 11536 17170 0 _024_
rlabel metal1 17112 12818 17112 12818 0 _025_
rlabel metal1 15977 16490 15977 16490 0 _026_
rlabel via1 17245 15402 17245 15402 0 _027_
rlabel metal1 14904 12410 14904 12410 0 _028_
rlabel metal1 13248 13158 13248 13158 0 _029_
rlabel metal3 18124 13532 18124 13532 0 _030_
rlabel metal1 14214 12614 14214 12614 0 _031_
rlabel metal1 18354 14416 18354 14416 0 _032_
rlabel metal2 17066 13770 17066 13770 0 _033_
rlabel metal1 13800 16150 13800 16150 0 _034_
rlabel metal1 16698 13294 16698 13294 0 _035_
rlabel metal1 17250 13362 17250 13362 0 _036_
rlabel metal1 17388 13498 17388 13498 0 _037_
rlabel metal1 16146 13770 16146 13770 0 _038_
rlabel metal1 7314 15538 7314 15538 0 _039_
rlabel metal1 8418 15436 8418 15436 0 _040_
rlabel metal1 9154 15470 9154 15470 0 _041_
rlabel metal2 10810 16660 10810 16660 0 _042_
rlabel metal1 10580 15062 10580 15062 0 _043_
rlabel viali 10349 14994 10349 14994 0 _044_
rlabel metal2 12834 15776 12834 15776 0 _045_
rlabel metal1 9568 14246 9568 14246 0 _046_
rlabel metal1 13064 14314 13064 14314 0 _047_
rlabel metal1 10212 14382 10212 14382 0 _048_
rlabel metal2 9522 15130 9522 15130 0 _049_
rlabel metal1 9844 14586 9844 14586 0 _050_
rlabel metal2 6578 16864 6578 16864 0 _051_
rlabel metal1 3818 15878 3818 15878 0 _052_
rlabel metal1 4370 16592 4370 16592 0 _053_
rlabel metal1 2530 15504 2530 15504 0 _054_
rlabel metal2 9890 14756 9890 14756 0 _055_
rlabel metal2 3818 15980 3818 15980 0 _056_
rlabel via1 4001 14994 4001 14994 0 _057_
rlabel metal2 4094 15504 4094 15504 0 _058_
rlabel metal1 4646 14858 4646 14858 0 _059_
rlabel metal1 4186 6834 4186 6834 0 _060_
rlabel metal2 5106 15300 5106 15300 0 _061_
rlabel metal1 6118 15572 6118 15572 0 _062_
rlabel metal1 2438 15470 2438 15470 0 _063_
rlabel metal2 1978 14246 1978 14246 0 _064_
rlabel metal2 2070 9316 2070 9316 0 _065_
rlabel metal1 1702 7854 1702 7854 0 _066_
rlabel metal1 1932 10506 1932 10506 0 _067_
rlabel metal1 4623 10030 4623 10030 0 _068_
rlabel metal2 4278 10778 4278 10778 0 _069_
rlabel metal1 4095 10064 4095 10064 0 _070_
rlabel metal2 4462 9690 4462 9690 0 _071_
rlabel metal1 4876 10234 4876 10234 0 _072_
rlabel metal2 3634 7684 3634 7684 0 _073_
rlabel metal1 5060 11118 5060 11118 0 _074_
rlabel metal1 4186 9418 4186 9418 0 _075_
rlabel metal1 2392 10574 2392 10574 0 _076_
rlabel metal1 1840 8534 1840 8534 0 _077_
rlabel metal1 2599 6766 2599 6766 0 _078_
rlabel metal1 1794 12172 1794 12172 0 _079_
rlabel metal1 4278 7480 4278 7480 0 _080_
rlabel metal1 2300 7378 2300 7378 0 _081_
rlabel metal2 2622 8415 2622 8415 0 _082_
rlabel metal1 1978 8296 1978 8296 0 _083_
rlabel metal1 2254 8602 2254 8602 0 _084_
rlabel metal1 4140 12614 4140 12614 0 _085_
rlabel metal1 5382 10234 5382 10234 0 _086_
rlabel metal2 1150 9044 1150 9044 0 _087_
rlabel metal1 3634 12784 3634 12784 0 _088_
rlabel metal1 3818 12648 3818 12648 0 _089_
rlabel metal1 1748 12954 1748 12954 0 _090_
rlabel metal2 5750 10574 5750 10574 0 _091_
rlabel metal1 4002 6630 4002 6630 0 _092_
rlabel via2 1150 11611 1150 11611 0 _093_
rlabel metal1 5014 8500 5014 8500 0 _094_
rlabel metal1 1932 13226 1932 13226 0 _095_
rlabel metal1 6348 12342 6348 12342 0 _096_
rlabel metal1 5382 7174 5382 7174 0 _097_
rlabel metal1 11638 12206 11638 12206 0 _098_
rlabel metal1 4462 14382 4462 14382 0 _099_
rlabel metal2 3910 14314 3910 14314 0 _100_
rlabel metal1 1656 14586 1656 14586 0 _101_
rlabel metal1 5152 14586 5152 14586 0 _102_
rlabel metal1 4784 12954 4784 12954 0 _103_
rlabel metal1 9384 10642 9384 10642 0 _104_
rlabel metal2 10442 12070 10442 12070 0 _105_
rlabel metal1 4324 13430 4324 13430 0 _106_
rlabel metal1 2392 13430 2392 13430 0 _107_
rlabel metal2 4554 13974 4554 13974 0 _108_
rlabel metal2 10902 12104 10902 12104 0 _109_
rlabel metal1 8004 13838 8004 13838 0 _110_
rlabel metal1 7084 13294 7084 13294 0 _111_
rlabel metal1 8280 15334 8280 15334 0 _112_
rlabel metal1 7958 14790 7958 14790 0 _113_
rlabel metal1 7084 14586 7084 14586 0 _114_
rlabel metal2 7774 13362 7774 13362 0 _115_
rlabel metal1 7498 14314 7498 14314 0 _116_
rlabel metal2 11178 16490 11178 16490 0 _117_
rlabel metal1 10672 12818 10672 12818 0 _118_
rlabel metal1 6854 15096 6854 15096 0 _119_
rlabel metal1 6992 14246 6992 14246 0 _120_
rlabel metal3 8211 16660 8211 16660 0 _121_
rlabel metal1 8188 13226 8188 13226 0 _122_
rlabel metal1 7406 14858 7406 14858 0 _123_
rlabel metal1 8832 11730 8832 11730 0 _124_
rlabel metal1 9062 13430 9062 13430 0 _125_
rlabel metal1 11316 14858 11316 14858 0 _126_
rlabel metal2 11178 13804 11178 13804 0 _127_
rlabel metal2 12788 13532 12788 13532 0 _128_
rlabel metal2 16974 13124 16974 13124 0 _129_
rlabel metal2 18078 13328 18078 13328 0 _130_
rlabel metal1 16560 11866 16560 11866 0 _131_
rlabel metal2 16422 11594 16422 11594 0 _132_
rlabel metal1 15426 13974 15426 13974 0 _133_
rlabel metal2 17894 14314 17894 14314 0 _134_
rlabel metal1 18354 15402 18354 15402 0 _135_
rlabel metal1 16836 13362 16836 13362 0 _136_
rlabel metal1 16882 14552 16882 14552 0 _137_
rlabel metal3 16054 14212 16054 14212 0 _138_
rlabel metal1 18446 13770 18446 13770 0 _139_
rlabel metal1 16146 13498 16146 13498 0 _140_
rlabel metal2 12926 13549 12926 13549 0 _141_
rlabel metal1 17618 12682 17618 12682 0 _142_
rlabel metal1 15489 12954 15489 12954 0 _143_
rlabel metal1 16974 12614 16974 12614 0 _144_
rlabel metal1 14444 12818 14444 12818 0 _145_
rlabel metal1 9752 12818 9752 12818 0 _146_
rlabel metal2 15042 16116 15042 16116 0 _147_
rlabel metal1 14306 16048 14306 16048 0 _148_
rlabel metal1 15732 15674 15732 15674 0 _149_
rlabel metal1 16192 14994 16192 14994 0 _150_
rlabel metal1 18078 14416 18078 14416 0 _151_
rlabel metal1 18538 13498 18538 13498 0 _152_
rlabel metal2 15686 13039 15686 13039 0 io_in[10]
rlabel metal3 18546 14484 18546 14484 0 io_in[11]
rlabel metal3 15479 12988 15479 12988 0 io_in[12]
rlabel metal1 15042 16694 15042 16694 0 io_in[13]
rlabel metal3 19236 18156 19236 18156 0 io_in[14]
rlabel metal2 19320 19244 19320 19244 0 io_in[15]
rlabel metal2 17526 19244 17526 19244 0 io_in[16]
rlabel metal1 14996 13294 14996 13294 0 io_in[17]
rlabel metal1 14490 15504 14490 15504 0 io_in[18]
rlabel metal2 13754 17340 13754 17340 0 io_in[19]
rlabel metal2 8464 14076 8464 14076 0 io_in[20]
rlabel metal2 6670 11662 6670 11662 0 io_in[21]
rlabel metal3 6532 12852 6532 12852 0 io_in[22]
rlabel metal2 1932 12988 1932 12988 0 io_in[23]
rlabel metal3 3419 18292 3419 18292 0 io_in[24]
rlabel metal2 7130 8160 7130 8160 0 io_in[25]
rlabel metal3 1717 15844 1717 15844 0 io_in[26]
rlabel metal3 1855 14620 1855 14620 0 io_in[27]
rlabel metal2 4370 8823 4370 8823 0 io_in[28]
rlabel metal1 5750 10642 5750 10642 0 io_in[29]
rlabel metal1 7682 11118 7682 11118 0 io_in[30]
rlabel metal1 5796 8466 5796 8466 0 io_in[31]
rlabel metal1 6762 8432 6762 8432 0 io_in[32]
rlabel metal1 4830 6732 4830 6732 0 io_in[33]
rlabel metal1 4370 6324 4370 6324 0 io_in[34]
rlabel metal2 17710 10897 17710 10897 0 io_in[8]
rlabel metal1 17296 9078 17296 9078 0 io_in[9]
rlabel metal3 1188 4420 1188 4420 0 io_out[35]
rlabel metal1 14766 14314 14766 14314 0 mod.clock_counter_a\[0\]
rlabel metal1 15180 14382 15180 14382 0 mod.clock_counter_a\[1\]
rlabel metal1 16054 14960 16054 14960 0 mod.clock_counter_a\[2\]
rlabel metal1 15778 15028 15778 15028 0 mod.clock_counter_a\[3\]
rlabel viali 15221 15470 15221 15470 0 mod.clock_counter_a\[4\]
rlabel metal1 17112 16558 17112 16558 0 mod.clock_counter_a\[5\]
rlabel metal2 18354 16388 18354 16388 0 mod.clock_counter_a\[6\]
rlabel metal1 13018 16014 13018 16014 0 mod.clock_counter_b\[0\]
rlabel metal1 7912 14586 7912 14586 0 mod.clock_counter_b\[1\]
rlabel metal1 12834 16116 12834 16116 0 mod.clock_counter_b\[2\]
rlabel metal1 10718 13940 10718 13940 0 mod.clock_counter_b\[3\]
rlabel metal2 12650 15232 12650 15232 0 mod.clock_counter_b\[4\]
rlabel metal1 13064 15402 13064 15402 0 mod.clock_counter_b\[5\]
rlabel metal1 12765 17306 12765 17306 0 mod.clock_counter_b\[6\]
rlabel metal1 6026 7310 6026 7310 0 mod.clock_counter_c\[0\]
rlabel metal1 5198 7446 5198 7446 0 mod.clock_counter_c\[1\]
rlabel metal1 5290 15334 5290 15334 0 mod.clock_counter_c\[2\]
rlabel metal1 3956 16558 3956 16558 0 mod.clock_counter_c\[3\]
rlabel metal1 5336 14790 5336 14790 0 mod.clock_counter_c\[4\]
rlabel metal1 5244 14314 5244 14314 0 mod.clock_counter_c\[5\]
rlabel metal2 1610 15946 1610 15946 0 mod.clock_counter_c\[6\]
rlabel metal1 3358 12682 3358 12682 0 mod.clock_counter_d\[0\]
rlabel metal2 2714 8228 2714 8228 0 mod.clock_counter_d\[1\]
rlabel metal1 4278 9962 4278 9962 0 mod.clock_counter_d\[2\]
rlabel metal1 5152 12138 5152 12138 0 mod.clock_counter_d\[3\]
rlabel metal1 6762 10608 6762 10608 0 mod.clock_counter_d\[4\]
rlabel metal1 3542 8500 3542 8500 0 mod.clock_counter_d\[5\]
rlabel metal1 3450 10608 3450 10608 0 mod.clock_counter_d\[6\]
rlabel metal1 6302 9996 6302 9996 0 mod.clock_syn
rlabel metal2 11270 13770 11270 13770 0 mod.div_clock\[0\]
rlabel metal1 9936 14042 9936 14042 0 mod.div_clock\[1\]
rlabel metal1 6854 13702 6854 13702 0 mod.div_clock\[2\]
rlabel metal1 7866 12954 7866 12954 0 mod.div_clock\[3\]
rlabel metal2 15502 12767 15502 12767 0 net1
rlabel metal1 13018 17000 13018 17000 0 net10
rlabel metal2 7314 11492 7314 11492 0 net100
rlabel metal2 4002 9299 4002 9299 0 net101
rlabel metal3 1027 9316 1027 9316 0 net102
rlabel metal1 2990 5882 2990 5882 0 net103
rlabel metal2 2806 6035 2806 6035 0 net104
rlabel via2 4002 5661 4002 5661 0 net105
rlabel metal2 1610 3111 1610 3111 0 net106
rlabel metal3 1464 1972 1464 1972 0 net107
rlabel metal2 13110 13401 13110 13401 0 net11
rlabel metal2 6854 11764 6854 11764 0 net12
rlabel metal1 8326 11322 8326 11322 0 net13
rlabel metal3 7291 16524 7291 16524 0 net14
rlabel metal1 5842 16014 5842 16014 0 net15
rlabel metal1 8188 8058 8188 8058 0 net16
rlabel metal1 4462 6766 4462 6766 0 net17
rlabel metal1 7222 9078 7222 9078 0 net18
rlabel metal1 6256 8602 6256 8602 0 net19
rlabel metal1 17526 13226 17526 13226 0 net2
rlabel metal2 2622 11594 2622 11594 0 net20
rlabel metal1 5106 11730 5106 11730 0 net21
rlabel metal1 4830 7888 4830 7888 0 net22
rlabel metal1 1794 5644 1794 5644 0 net23
rlabel metal1 1794 5236 1794 5236 0 net24
rlabel metal1 3956 6290 3956 6290 0 net25
rlabel metal1 17434 11322 17434 11322 0 net26
rlabel metal1 15732 10982 15732 10982 0 net27
rlabel metal2 6118 7242 6118 7242 0 net28
rlabel metal1 1610 9588 1610 9588 0 net29
rlabel metal1 15686 14382 15686 14382 0 net3
rlabel metal1 1656 16082 1656 16082 0 net30
rlabel metal2 8602 17374 8602 17374 0 net31
rlabel metal1 11224 14994 11224 14994 0 net32
rlabel metal2 18354 2125 18354 2125 0 net33
rlabel metal2 18354 3281 18354 3281 0 net34
rlabel metal1 18768 4590 18768 4590 0 net35
rlabel via2 18354 5661 18354 5661 0 net36
rlabel via2 18354 6749 18354 6749 0 net37
rlabel via2 18354 7939 18354 7939 0 net38
rlabel via2 18354 9163 18354 9163 0 net39
rlabel metal1 14858 12648 14858 12648 0 net4
rlabel metal2 18354 10319 18354 10319 0 net40
rlabel via2 17526 11611 17526 11611 0 net41
rlabel metal3 18178 12852 18178 12852 0 net42
rlabel metal1 14214 13838 14214 13838 0 net43
rlabel metal1 13662 13362 13662 13362 0 net44
rlabel metal2 14260 13804 14260 13804 0 net45
rlabel via3 16261 12444 16261 12444 0 net46
rlabel metal3 15847 13124 15847 13124 0 net47
rlabel metal1 18676 15878 18676 15878 0 net48
rlabel metal1 13570 13906 13570 13906 0 net49
rlabel metal1 14168 12750 14168 12750 0 net5
rlabel metal1 14076 14586 14076 14586 0 net50
rlabel metal2 14306 16762 14306 16762 0 net51
rlabel metal2 9246 17452 9246 17452 0 net52
rlabel metal1 7084 11730 7084 11730 0 net53
rlabel metal3 5037 15980 5037 15980 0 net54
rlabel metal2 2622 16585 2622 16585 0 net55
rlabel metal2 414 18897 414 18897 0 net56
rlabel metal3 1717 17476 1717 17476 0 net57
rlabel metal3 2499 16252 2499 16252 0 net58
rlabel metal3 1786 15028 1786 15028 0 net59
rlabel metal1 15778 9418 15778 9418 0 net6
rlabel metal1 7682 10574 7682 10574 0 net60
rlabel metal3 1740 12580 1740 12580 0 net61
rlabel metal2 6762 10642 6762 10642 0 net62
rlabel metal3 1717 10132 1717 10132 0 net63
rlabel metal1 3220 6290 3220 6290 0 net64
rlabel metal1 4554 7310 4554 7310 0 net65
rlabel metal2 2898 5831 2898 5831 0 net66
rlabel metal2 1610 4675 1610 4675 0 net67
rlabel metal2 1610 3859 1610 3859 0 net68
rlabel metal3 1142 2788 1142 2788 0 net69
rlabel metal2 17434 10642 17434 10642 0 net7
rlabel metal3 1786 1564 1786 1564 0 net70
rlabel metal2 17710 1921 17710 1921 0 net71
rlabel metal3 18868 2652 18868 2652 0 net72
rlabel via2 18354 3893 18354 3893 0 net73
rlabel via2 18354 5083 18354 5083 0 net74
rlabel via2 18354 6307 18354 6307 0 net75
rlabel via2 18354 7395 18354 7395 0 net76
rlabel metal1 18768 8466 18768 8466 0 net77
rlabel metal2 18354 9775 18354 9775 0 net78
rlabel metal2 18354 10931 18354 10931 0 net79
rlabel metal2 11914 14756 11914 14756 0 net8
rlabel via2 16330 12699 16330 12699 0 net80
rlabel metal3 16905 13396 16905 13396 0 net81
rlabel metal2 16008 13668 16008 13668 0 net82
rlabel metal2 18722 12444 18722 12444 0 net83
rlabel metal2 14490 11305 14490 11305 0 net84
rlabel metal3 16545 18564 16545 18564 0 net85
rlabel metal1 19136 17510 19136 17510 0 net86
rlabel metal1 14996 12818 14996 12818 0 net87
rlabel metal1 14352 13906 14352 13906 0 net88
rlabel metal1 12282 14994 12282 14994 0 net89
rlabel metal2 13294 16082 13294 16082 0 net9
rlabel metal2 13570 16660 13570 16660 0 net90
rlabel metal2 7866 17068 7866 17068 0 net91
rlabel metal2 7406 11492 7406 11492 0 net92
rlabel metal3 5957 16116 5957 16116 0 net93
rlabel metal2 828 19244 828 19244 0 net94
rlabel metal3 4983 17884 4983 17884 0 net95
rlabel metal3 5842 16864 5842 16864 0 net96
rlabel metal3 1832 15436 1832 15436 0 net97
rlabel metal3 2154 14212 2154 14212 0 net98
rlabel metal2 11546 13396 11546 13396 0 net99
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
