magic
tech sky130A
magscale 1 2
timestamp 1672340475
<< obsli1 >>
rect 1104 2159 22816 27761
<< obsm1 >>
rect 1104 2128 22976 27872
<< metal2 >>
rect 1214 29200 1270 30000
rect 2042 29200 2098 30000
rect 2870 29200 2926 30000
rect 3698 29200 3754 30000
rect 4526 29200 4582 30000
rect 5354 29200 5410 30000
rect 6182 29200 6238 30000
rect 7010 29200 7066 30000
rect 7838 29200 7894 30000
rect 8666 29200 8722 30000
rect 9494 29200 9550 30000
rect 10322 29200 10378 30000
rect 11150 29200 11206 30000
rect 11978 29200 12034 30000
rect 12806 29200 12862 30000
rect 13634 29200 13690 30000
rect 14462 29200 14518 30000
rect 15290 29200 15346 30000
rect 16118 29200 16174 30000
rect 16946 29200 17002 30000
rect 17774 29200 17830 30000
rect 18602 29200 18658 30000
rect 19430 29200 19486 30000
rect 20258 29200 20314 30000
rect 21086 29200 21142 30000
rect 21914 29200 21970 30000
rect 22742 29200 22798 30000
<< obsm2 >>
rect 1326 29144 1986 29322
rect 2154 29144 2814 29322
rect 2982 29144 3642 29322
rect 3810 29144 4470 29322
rect 4638 29144 5298 29322
rect 5466 29144 6126 29322
rect 6294 29144 6954 29322
rect 7122 29144 7782 29322
rect 7950 29144 8610 29322
rect 8778 29144 9438 29322
rect 9606 29144 10266 29322
rect 10434 29144 11094 29322
rect 11262 29144 11922 29322
rect 12090 29144 12750 29322
rect 12918 29144 13578 29322
rect 13746 29144 14406 29322
rect 14574 29144 15234 29322
rect 15402 29144 16062 29322
rect 16230 29144 16890 29322
rect 17058 29144 17718 29322
rect 17886 29144 18546 29322
rect 18714 29144 19374 29322
rect 19542 29144 20202 29322
rect 20370 29144 21030 29322
rect 21198 29144 21858 29322
rect 22026 29144 22686 29322
rect 22854 29144 22970 29322
rect 1214 983 22970 29144
<< metal3 >>
rect 0 28840 800 28960
rect 0 28160 800 28280
rect 0 27480 800 27600
rect 0 26800 800 26920
rect 23200 26800 24000 26920
rect 0 26120 800 26240
rect 23200 26256 24000 26376
rect 23200 25712 24000 25832
rect 0 25440 800 25560
rect 23200 25168 24000 25288
rect 0 24760 800 24880
rect 23200 24624 24000 24744
rect 0 24080 800 24200
rect 23200 24080 24000 24200
rect 0 23400 800 23520
rect 23200 23536 24000 23656
rect 23200 22992 24000 23112
rect 0 22720 800 22840
rect 23200 22448 24000 22568
rect 0 22040 800 22160
rect 23200 21904 24000 22024
rect 0 21360 800 21480
rect 23200 21360 24000 21480
rect 0 20680 800 20800
rect 23200 20816 24000 20936
rect 23200 20272 24000 20392
rect 0 20000 800 20120
rect 23200 19728 24000 19848
rect 0 19320 800 19440
rect 23200 19184 24000 19304
rect 0 18640 800 18760
rect 23200 18640 24000 18760
rect 0 17960 800 18080
rect 23200 18096 24000 18216
rect 23200 17552 24000 17672
rect 0 17280 800 17400
rect 23200 17008 24000 17128
rect 0 16600 800 16720
rect 23200 16464 24000 16584
rect 0 15920 800 16040
rect 23200 15920 24000 16040
rect 0 15240 800 15360
rect 23200 15376 24000 15496
rect 23200 14832 24000 14952
rect 0 14560 800 14680
rect 23200 14288 24000 14408
rect 0 13880 800 14000
rect 23200 13744 24000 13864
rect 0 13200 800 13320
rect 23200 13200 24000 13320
rect 0 12520 800 12640
rect 23200 12656 24000 12776
rect 23200 12112 24000 12232
rect 0 11840 800 11960
rect 23200 11568 24000 11688
rect 0 11160 800 11280
rect 23200 11024 24000 11144
rect 0 10480 800 10600
rect 23200 10480 24000 10600
rect 0 9800 800 9920
rect 23200 9936 24000 10056
rect 23200 9392 24000 9512
rect 0 9120 800 9240
rect 23200 8848 24000 8968
rect 0 8440 800 8560
rect 23200 8304 24000 8424
rect 0 7760 800 7880
rect 23200 7760 24000 7880
rect 0 7080 800 7200
rect 23200 7216 24000 7336
rect 23200 6672 24000 6792
rect 0 6400 800 6520
rect 23200 6128 24000 6248
rect 0 5720 800 5840
rect 23200 5584 24000 5704
rect 0 5040 800 5160
rect 23200 5040 24000 5160
rect 0 4360 800 4480
rect 23200 4496 24000 4616
rect 23200 3952 24000 4072
rect 0 3680 800 3800
rect 23200 3408 24000 3528
rect 0 3000 800 3120
rect 23200 2864 24000 2984
rect 0 2320 800 2440
rect 0 1640 800 1760
rect 0 960 800 1080
<< obsm3 >>
rect 880 28760 23200 28933
rect 800 28360 23200 28760
rect 880 28080 23200 28360
rect 800 27680 23200 28080
rect 880 27400 23200 27680
rect 800 27000 23200 27400
rect 880 26720 23120 27000
rect 800 26456 23200 26720
rect 800 26320 23120 26456
rect 880 26176 23120 26320
rect 880 26040 23200 26176
rect 800 25912 23200 26040
rect 800 25640 23120 25912
rect 880 25632 23120 25640
rect 880 25368 23200 25632
rect 880 25360 23120 25368
rect 800 25088 23120 25360
rect 800 24960 23200 25088
rect 880 24824 23200 24960
rect 880 24680 23120 24824
rect 800 24544 23120 24680
rect 800 24280 23200 24544
rect 880 24000 23120 24280
rect 800 23736 23200 24000
rect 800 23600 23120 23736
rect 880 23456 23120 23600
rect 880 23320 23200 23456
rect 800 23192 23200 23320
rect 800 22920 23120 23192
rect 880 22912 23120 22920
rect 880 22648 23200 22912
rect 880 22640 23120 22648
rect 800 22368 23120 22640
rect 800 22240 23200 22368
rect 880 22104 23200 22240
rect 880 21960 23120 22104
rect 800 21824 23120 21960
rect 800 21560 23200 21824
rect 880 21280 23120 21560
rect 800 21016 23200 21280
rect 800 20880 23120 21016
rect 880 20736 23120 20880
rect 880 20600 23200 20736
rect 800 20472 23200 20600
rect 800 20200 23120 20472
rect 880 20192 23120 20200
rect 880 19928 23200 20192
rect 880 19920 23120 19928
rect 800 19648 23120 19920
rect 800 19520 23200 19648
rect 880 19384 23200 19520
rect 880 19240 23120 19384
rect 800 19104 23120 19240
rect 800 18840 23200 19104
rect 880 18560 23120 18840
rect 800 18296 23200 18560
rect 800 18160 23120 18296
rect 880 18016 23120 18160
rect 880 17880 23200 18016
rect 800 17752 23200 17880
rect 800 17480 23120 17752
rect 880 17472 23120 17480
rect 880 17208 23200 17472
rect 880 17200 23120 17208
rect 800 16928 23120 17200
rect 800 16800 23200 16928
rect 880 16664 23200 16800
rect 880 16520 23120 16664
rect 800 16384 23120 16520
rect 800 16120 23200 16384
rect 880 15840 23120 16120
rect 800 15576 23200 15840
rect 800 15440 23120 15576
rect 880 15296 23120 15440
rect 880 15160 23200 15296
rect 800 15032 23200 15160
rect 800 14760 23120 15032
rect 880 14752 23120 14760
rect 880 14488 23200 14752
rect 880 14480 23120 14488
rect 800 14208 23120 14480
rect 800 14080 23200 14208
rect 880 13944 23200 14080
rect 880 13800 23120 13944
rect 800 13664 23120 13800
rect 800 13400 23200 13664
rect 880 13120 23120 13400
rect 800 12856 23200 13120
rect 800 12720 23120 12856
rect 880 12576 23120 12720
rect 880 12440 23200 12576
rect 800 12312 23200 12440
rect 800 12040 23120 12312
rect 880 12032 23120 12040
rect 880 11768 23200 12032
rect 880 11760 23120 11768
rect 800 11488 23120 11760
rect 800 11360 23200 11488
rect 880 11224 23200 11360
rect 880 11080 23120 11224
rect 800 10944 23120 11080
rect 800 10680 23200 10944
rect 880 10400 23120 10680
rect 800 10136 23200 10400
rect 800 10000 23120 10136
rect 880 9856 23120 10000
rect 880 9720 23200 9856
rect 800 9592 23200 9720
rect 800 9320 23120 9592
rect 880 9312 23120 9320
rect 880 9048 23200 9312
rect 880 9040 23120 9048
rect 800 8768 23120 9040
rect 800 8640 23200 8768
rect 880 8504 23200 8640
rect 880 8360 23120 8504
rect 800 8224 23120 8360
rect 800 7960 23200 8224
rect 880 7680 23120 7960
rect 800 7416 23200 7680
rect 800 7280 23120 7416
rect 880 7136 23120 7280
rect 880 7000 23200 7136
rect 800 6872 23200 7000
rect 800 6600 23120 6872
rect 880 6592 23120 6600
rect 880 6328 23200 6592
rect 880 6320 23120 6328
rect 800 6048 23120 6320
rect 800 5920 23200 6048
rect 880 5784 23200 5920
rect 880 5640 23120 5784
rect 800 5504 23120 5640
rect 800 5240 23200 5504
rect 880 4960 23120 5240
rect 800 4696 23200 4960
rect 800 4560 23120 4696
rect 880 4416 23120 4560
rect 880 4280 23200 4416
rect 800 4152 23200 4280
rect 800 3880 23120 4152
rect 880 3872 23120 3880
rect 880 3608 23200 3872
rect 880 3600 23120 3608
rect 800 3328 23120 3600
rect 800 3200 23200 3328
rect 880 3064 23200 3200
rect 880 2920 23120 3064
rect 800 2784 23120 2920
rect 800 2520 23200 2784
rect 880 2240 23200 2520
rect 800 1840 23200 2240
rect 880 1560 23200 1840
rect 800 1160 23200 1560
rect 880 987 23200 1160
<< metal4 >>
rect 3658 2128 3978 27792
rect 6372 2128 6692 27792
rect 9086 2128 9406 27792
rect 11800 2128 12120 27792
rect 14514 2128 14834 27792
rect 17228 2128 17548 27792
rect 19942 2128 20262 27792
rect 22656 2128 22976 27792
<< obsm4 >>
rect 4107 14451 6292 26485
rect 6772 14451 9006 26485
rect 9486 14451 11720 26485
rect 12200 14451 14434 26485
rect 14914 14451 17148 26485
rect 17628 14451 19862 26485
rect 20342 14451 21469 26485
<< labels >>
rlabel metal3 s 23200 2864 24000 2984 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 23200 19184 24000 19304 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 23200 20816 24000 20936 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 23200 22448 24000 22568 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 23200 24080 24000 24200 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 23200 25712 24000 25832 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 22742 29200 22798 30000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 20258 29200 20314 30000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 17774 29200 17830 30000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 15290 29200 15346 30000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 12806 29200 12862 30000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 23200 4496 24000 4616 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 10322 29200 10378 30000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 7838 29200 7894 30000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 5354 29200 5410 30000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 2870 29200 2926 30000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 23200 6128 24000 6248 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 23200 7760 24000 7880 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 23200 9392 24000 9512 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 23200 11024 24000 11144 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 23200 12656 24000 12776 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 23200 14288 24000 14408 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 23200 15920 24000 16040 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 23200 17552 24000 17672 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 23200 3952 24000 4072 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 23200 20272 24000 20392 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 23200 21904 24000 22024 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 23200 23536 24000 23656 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 23200 25168 24000 25288 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 23200 26800 24000 26920 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 21086 29200 21142 30000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 18602 29200 18658 30000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 13634 29200 13690 30000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 11150 29200 11206 30000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 23200 5584 24000 5704 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 8666 29200 8722 30000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 6182 29200 6238 30000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 3698 29200 3754 30000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 1214 29200 1270 30000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 23200 7216 24000 7336 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 960 800 1080 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 23200 8848 24000 8968 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 23200 10480 24000 10600 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 23200 12112 24000 12232 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 23200 13744 24000 13864 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 23200 15376 24000 15496 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 23200 17008 24000 17128 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 23200 18640 24000 18760 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 23200 3408 24000 3528 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 23200 19728 24000 19848 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 23200 21360 24000 21480 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 23200 22992 24000 23112 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 23200 24624 24000 24744 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 23200 26256 24000 26376 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 21914 29200 21970 30000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 19430 29200 19486 30000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 16946 29200 17002 30000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 14462 29200 14518 30000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 11978 29200 12034 30000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 23200 5040 24000 5160 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 9494 29200 9550 30000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 7010 29200 7066 30000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 4526 29200 4582 30000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 2042 29200 2098 30000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 23200 6672 24000 6792 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 23200 8304 24000 8424 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 23200 9936 24000 10056 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 23200 11568 24000 11688 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 23200 13200 24000 13320 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 23200 14832 24000 14952 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 23200 16464 24000 16584 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 23200 18096 24000 18216 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 3658 2128 3978 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 9086 2128 9406 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 14514 2128 14834 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19942 2128 20262 27792 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 11800 2128 12120 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 17228 2128 17548 27792 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 22656 2128 22976 27792 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1085150
string GDS_FILE /home/runner/work/clock_divide_select_4ch_tiny_user/clock_divide_select_4ch_tiny_user/openlane/tiny_user_project/runs/22_12_29_18_59/results/signoff/tiny_user_project.magic.gds
string GDS_START 153314
<< end >>

