magic
tech sky130A
magscale 1 2
timestamp 1672340473
<< viali >>
rect 9321 27625 9355 27659
rect 4721 27557 4755 27591
rect 8585 27557 8619 27591
rect 15485 27557 15519 27591
rect 17509 27557 17543 27591
rect 20085 27557 20119 27591
rect 20729 27557 20763 27591
rect 7205 27489 7239 27523
rect 12725 27489 12759 27523
rect 15393 27489 15427 27523
rect 18797 27489 18831 27523
rect 1593 27421 1627 27455
rect 2237 27421 2271 27455
rect 3065 27421 3099 27455
rect 5181 27421 5215 27455
rect 5365 27421 5399 27455
rect 5825 27421 5859 27455
rect 6561 27421 6595 27455
rect 6745 27421 6779 27455
rect 11161 27421 11195 27455
rect 11713 27421 11747 27455
rect 12541 27421 12575 27455
rect 12909 27421 12943 27455
rect 13093 27421 13127 27455
rect 14468 27421 14502 27455
rect 14565 27421 14599 27455
rect 14785 27421 14819 27455
rect 14933 27421 14967 27455
rect 17049 27421 17083 27455
rect 18337 27421 18371 27455
rect 19441 27421 19475 27455
rect 21281 27421 21315 27455
rect 22109 27421 22143 27455
rect 7450 27353 7484 27387
rect 10894 27353 10928 27387
rect 14657 27353 14691 27387
rect 15853 27353 15887 27387
rect 1777 27285 1811 27319
rect 2421 27285 2455 27319
rect 2973 27285 3007 27319
rect 4077 27285 4111 27319
rect 5365 27285 5399 27319
rect 6009 27285 6043 27319
rect 6745 27285 6779 27319
rect 9781 27285 9815 27319
rect 11805 27285 11839 27319
rect 14289 27285 14323 27319
rect 16865 27285 16899 27319
rect 18153 27285 18187 27319
rect 21373 27285 21407 27319
rect 22201 27285 22235 27319
rect 7179 27081 7213 27115
rect 7941 27081 7975 27115
rect 14105 27081 14139 27115
rect 14565 27081 14599 27115
rect 20545 27081 20579 27115
rect 1593 27013 1627 27047
rect 1809 27013 1843 27047
rect 7389 27013 7423 27047
rect 9137 27013 9171 27047
rect 15025 27013 15059 27047
rect 2421 26945 2455 26979
rect 3801 26945 3835 26979
rect 4537 26945 4571 26979
rect 5181 26945 5215 26979
rect 5825 26945 5859 26979
rect 7849 26945 7883 26979
rect 8125 26945 8159 26979
rect 10894 26945 10928 26979
rect 12837 26945 12871 26979
rect 13553 26945 13587 26979
rect 13829 26945 13863 26979
rect 13921 26945 13955 26979
rect 15577 26945 15611 26979
rect 16865 26945 16899 26979
rect 17785 26945 17819 26979
rect 19257 26945 19291 26979
rect 20361 26945 20395 26979
rect 22201 26945 22235 26979
rect 11161 26877 11195 26911
rect 13093 26877 13127 26911
rect 18613 26877 18647 26911
rect 6009 26809 6043 26843
rect 8769 26809 8803 26843
rect 14749 26809 14783 26843
rect 15761 26809 15795 26843
rect 16221 26809 16255 26843
rect 19901 26809 19935 26843
rect 1777 26741 1811 26775
rect 1961 26741 1995 26775
rect 2605 26741 2639 26775
rect 3065 26741 3099 26775
rect 5365 26741 5399 26775
rect 7021 26741 7055 26775
rect 7205 26741 7239 26775
rect 8309 26741 8343 26775
rect 9137 26741 9171 26775
rect 9321 26741 9355 26775
rect 9781 26741 9815 26775
rect 11713 26741 11747 26775
rect 13645 26741 13679 26775
rect 17969 26741 18003 26775
rect 21465 26741 21499 26775
rect 22017 26741 22051 26775
rect 2053 26537 2087 26571
rect 6929 26537 6963 26571
rect 7389 26537 7423 26571
rect 8401 26537 8435 26571
rect 8585 26537 8619 26571
rect 10057 26537 10091 26571
rect 10241 26537 10275 26571
rect 14473 26537 14507 26571
rect 1961 26469 1995 26503
rect 2789 26469 2823 26503
rect 4629 26469 4663 26503
rect 5641 26469 5675 26503
rect 12081 26469 12115 26503
rect 14289 26469 14323 26503
rect 15117 26469 15151 26503
rect 2513 26401 2547 26435
rect 6285 26401 6319 26435
rect 21649 26401 21683 26435
rect 3985 26333 4019 26367
rect 4813 26333 4847 26367
rect 5457 26333 5491 26367
rect 6745 26333 6779 26367
rect 7757 26333 7791 26367
rect 9689 26333 9723 26367
rect 10701 26333 10735 26367
rect 12541 26333 12575 26367
rect 12817 26333 12851 26367
rect 12909 26333 12943 26367
rect 13737 26333 13771 26367
rect 15945 26333 15979 26367
rect 16405 26333 16439 26367
rect 18889 26333 18923 26367
rect 19533 26333 19567 26367
rect 20361 26333 20395 26367
rect 1593 26265 1627 26299
rect 4077 26265 4111 26299
rect 7573 26265 7607 26299
rect 8217 26265 8251 26299
rect 8417 26265 8451 26299
rect 9229 26265 9263 26299
rect 10946 26265 10980 26299
rect 12725 26265 12759 26299
rect 14441 26265 14475 26299
rect 14657 26265 14691 26299
rect 18153 26265 18187 26299
rect 19625 26265 19659 26299
rect 20821 26265 20855 26299
rect 21005 26265 21039 26299
rect 21189 26265 21223 26299
rect 21833 26265 21867 26299
rect 22017 26265 22051 26299
rect 2973 26197 3007 26231
rect 10057 26197 10091 26231
rect 13093 26197 13127 26231
rect 13553 26197 13587 26231
rect 15761 26197 15795 26231
rect 2697 25993 2731 26027
rect 11161 25993 11195 26027
rect 13185 25993 13219 26027
rect 1961 25925 1995 25959
rect 3709 25925 3743 25959
rect 9121 25925 9155 25959
rect 9321 25925 9355 25959
rect 2605 25857 2639 25891
rect 2881 25857 2915 25891
rect 3893 25857 3927 25891
rect 4353 25857 4387 25891
rect 4537 25857 4571 25891
rect 6561 25857 6595 25891
rect 7481 25857 7515 25891
rect 8309 25857 8343 25891
rect 9788 25857 9822 25891
rect 10037 25857 10071 25891
rect 11713 25857 11747 25891
rect 11989 25857 12023 25891
rect 12081 25857 12115 25891
rect 12725 25857 12759 25891
rect 13829 25857 13863 25891
rect 14013 25857 14047 25891
rect 18705 25857 18739 25891
rect 19165 25857 19199 25891
rect 19809 25857 19843 25891
rect 20453 25857 20487 25891
rect 21281 25857 21315 25891
rect 22017 25857 22051 25891
rect 5641 25789 5675 25823
rect 8125 25789 8159 25823
rect 14473 25789 14507 25823
rect 21097 25789 21131 25823
rect 1593 25721 1627 25755
rect 2145 25721 2179 25755
rect 4997 25721 5031 25755
rect 8953 25721 8987 25755
rect 13645 25721 13679 25755
rect 19349 25721 19383 25755
rect 1961 25653 1995 25687
rect 3065 25653 3099 25687
rect 3525 25653 3559 25687
rect 4445 25653 4479 25687
rect 7665 25653 7699 25687
rect 8493 25653 8527 25687
rect 9137 25653 9171 25687
rect 11805 25653 11839 25687
rect 12265 25653 12299 25687
rect 13001 25653 13035 25687
rect 15209 25653 15243 25687
rect 19993 25653 20027 25687
rect 20637 25653 20671 25687
rect 21465 25653 21499 25687
rect 22201 25653 22235 25687
rect 1593 25449 1627 25483
rect 6193 25449 6227 25483
rect 6837 25449 6871 25483
rect 7849 25449 7883 25483
rect 8493 25449 8527 25483
rect 13277 25449 13311 25483
rect 20085 25449 20119 25483
rect 20269 25449 20303 25483
rect 20913 25449 20947 25483
rect 4261 25381 4295 25415
rect 5549 25313 5583 25347
rect 2706 25245 2740 25279
rect 2973 25245 3007 25279
rect 5089 25245 5123 25279
rect 7021 25245 7055 25279
rect 7757 25245 7791 25279
rect 8401 25245 8435 25279
rect 9597 25245 9631 25279
rect 10425 25245 10459 25279
rect 10681 25245 10715 25279
rect 12265 25245 12299 25279
rect 12541 25245 12575 25279
rect 12725 25245 12759 25279
rect 13369 25245 13403 25279
rect 19441 25245 19475 25279
rect 22026 25245 22060 25279
rect 22293 25245 22327 25279
rect 3985 25177 4019 25211
rect 9781 25177 9815 25211
rect 12357 25177 12391 25211
rect 20453 25177 20487 25211
rect 4445 25109 4479 25143
rect 4905 25109 4939 25143
rect 9965 25109 9999 25143
rect 11805 25109 11839 25143
rect 17785 25109 17819 25143
rect 18245 25109 18279 25143
rect 18797 25109 18831 25143
rect 19625 25109 19659 25143
rect 20253 25109 20287 25143
rect 9939 24905 9973 24939
rect 12633 24905 12667 24939
rect 20085 24905 20119 24939
rect 3709 24837 3743 24871
rect 10149 24837 10183 24871
rect 10793 24837 10827 24871
rect 19449 24837 19483 24871
rect 2706 24769 2740 24803
rect 2973 24769 3007 24803
rect 3593 24769 3627 24803
rect 3801 24769 3835 24803
rect 3985 24769 4019 24803
rect 4905 24769 4939 24803
rect 5549 24769 5583 24803
rect 6561 24769 6595 24803
rect 7389 24769 7423 24803
rect 7849 24769 7883 24803
rect 8493 24769 8527 24803
rect 9137 24769 9171 24803
rect 11161 24769 11195 24803
rect 11713 24769 11747 24803
rect 12817 24769 12851 24803
rect 18613 24769 18647 24803
rect 19257 24769 19291 24803
rect 21209 24769 21243 24803
rect 22201 24769 22235 24803
rect 12173 24701 12207 24735
rect 21465 24701 21499 24735
rect 5365 24633 5399 24667
rect 9321 24633 9355 24667
rect 9781 24633 9815 24667
rect 10609 24633 10643 24667
rect 11989 24633 12023 24667
rect 18153 24633 18187 24667
rect 1593 24565 1627 24599
rect 3433 24565 3467 24599
rect 4445 24565 4479 24599
rect 4629 24565 4663 24599
rect 7205 24565 7239 24599
rect 8585 24565 8619 24599
rect 9965 24565 9999 24599
rect 10793 24565 10827 24599
rect 17509 24565 17543 24599
rect 18705 24565 18739 24599
rect 19625 24565 19659 24599
rect 22017 24565 22051 24599
rect 5181 24361 5215 24395
rect 8493 24361 8527 24395
rect 9597 24361 9631 24395
rect 10425 24361 10459 24395
rect 11713 24361 11747 24395
rect 17417 24361 17451 24395
rect 18705 24361 18739 24395
rect 18889 24361 18923 24395
rect 20085 24361 20119 24395
rect 20913 24361 20947 24395
rect 4997 24293 5031 24327
rect 6653 24293 6687 24327
rect 7297 24293 7331 24327
rect 7941 24293 7975 24327
rect 20453 24293 20487 24327
rect 4445 24225 4479 24259
rect 10885 24225 10919 24259
rect 12449 24225 12483 24259
rect 2706 24157 2740 24191
rect 2973 24157 3007 24191
rect 4169 24157 4203 24191
rect 4261 24157 4295 24191
rect 4537 24157 4571 24191
rect 6837 24157 6871 24191
rect 10241 24157 10275 24191
rect 11253 24157 11287 24191
rect 16773 24157 16807 24191
rect 17233 24157 17267 24191
rect 17877 24157 17911 24191
rect 18061 24157 18095 24191
rect 22026 24157 22060 24191
rect 22293 24157 22327 24191
rect 5365 24089 5399 24123
rect 6010 24089 6044 24123
rect 6193 24089 6227 24123
rect 11069 24089 11103 24123
rect 18521 24089 18555 24123
rect 1593 24021 1627 24055
rect 3985 24021 4019 24055
rect 5165 24021 5199 24055
rect 5825 24021 5859 24055
rect 18061 24021 18095 24055
rect 18721 24021 18755 24055
rect 19901 24021 19935 24055
rect 20085 24021 20119 24055
rect 3893 23817 3927 23851
rect 5825 23817 5859 23851
rect 6561 23817 6595 23851
rect 10977 23817 11011 23851
rect 17601 23817 17635 23851
rect 22017 23817 22051 23851
rect 8125 23749 8159 23783
rect 17417 23749 17451 23783
rect 18337 23749 18371 23783
rect 21220 23749 21254 23783
rect 1593 23681 1627 23715
rect 2145 23681 2179 23715
rect 2513 23681 2547 23715
rect 3065 23681 3099 23715
rect 3433 23681 3467 23715
rect 5006 23681 5040 23715
rect 5917 23681 5951 23715
rect 6745 23681 6779 23715
rect 6837 23681 6871 23715
rect 7389 23681 7423 23715
rect 7573 23681 7607 23715
rect 11161 23681 11195 23715
rect 17233 23681 17267 23715
rect 18061 23681 18095 23715
rect 18245 23681 18279 23715
rect 18429 23681 18463 23715
rect 19073 23681 19107 23715
rect 19349 23681 19383 23715
rect 19441 23681 19475 23715
rect 22201 23681 22235 23715
rect 2605 23613 2639 23647
rect 5273 23613 5307 23647
rect 19165 23613 19199 23647
rect 21465 23613 21499 23647
rect 19625 23545 19659 23579
rect 7481 23477 7515 23511
rect 18613 23477 18647 23511
rect 20085 23477 20119 23511
rect 2973 23273 3007 23307
rect 5917 23273 5951 23307
rect 7757 23273 7791 23307
rect 16865 23273 16899 23307
rect 19809 23273 19843 23307
rect 19993 23273 20027 23307
rect 7205 23205 7239 23239
rect 17049 23205 17083 23239
rect 17877 23205 17911 23239
rect 18705 23205 18739 23239
rect 18889 23205 18923 23239
rect 18429 23137 18463 23171
rect 21189 23137 21223 23171
rect 21649 23137 21683 23171
rect 1593 23069 1627 23103
rect 1860 23069 1894 23103
rect 4164 23069 4198 23103
rect 4353 23069 4387 23103
rect 4481 23069 4515 23103
rect 4629 23069 4663 23103
rect 5273 23069 5307 23103
rect 6101 23069 6135 23103
rect 6745 23069 6779 23103
rect 19441 23069 19475 23103
rect 20453 23069 20487 23103
rect 21281 23069 21315 23103
rect 21925 23069 21959 23103
rect 4261 23001 4295 23035
rect 5457 23001 5491 23035
rect 16681 23001 16715 23035
rect 16897 23001 16931 23035
rect 17509 23001 17543 23035
rect 3985 22933 4019 22967
rect 5089 22933 5123 22967
rect 6561 22933 6595 22967
rect 17969 22933 18003 22967
rect 19809 22933 19843 22967
rect 20729 22933 20763 22967
rect 7113 22729 7147 22763
rect 18245 22729 18279 22763
rect 18613 22729 18647 22763
rect 20085 22729 20119 22763
rect 22109 22729 22143 22763
rect 1860 22661 1894 22695
rect 3801 22661 3835 22695
rect 4445 22661 4479 22695
rect 4661 22661 4695 22695
rect 21220 22661 21254 22695
rect 1593 22593 1627 22627
rect 5917 22593 5951 22627
rect 6653 22593 6687 22627
rect 17509 22593 17543 22627
rect 17693 22593 17727 22627
rect 18153 22593 18187 22627
rect 18429 22593 18463 22627
rect 19257 22593 19291 22627
rect 19349 22593 19383 22627
rect 19625 22593 19659 22627
rect 22293 22593 22327 22627
rect 3433 22525 3467 22559
rect 19533 22525 19567 22559
rect 21465 22525 21499 22559
rect 2973 22457 3007 22491
rect 5273 22457 5307 22491
rect 3801 22389 3835 22423
rect 3985 22389 4019 22423
rect 4629 22389 4663 22423
rect 4813 22389 4847 22423
rect 17601 22389 17635 22423
rect 19073 22389 19107 22423
rect 4169 22185 4203 22219
rect 5457 22185 5491 22219
rect 20269 22185 20303 22219
rect 4353 22117 4387 22151
rect 1593 22049 1627 22083
rect 4905 22049 4939 22083
rect 6101 22049 6135 22083
rect 10609 22049 10643 22083
rect 18429 22049 18463 22083
rect 1860 21981 1894 22015
rect 4813 21981 4847 22015
rect 6561 21981 6595 22015
rect 10701 21981 10735 22015
rect 18613 21981 18647 22015
rect 18889 21981 18923 22015
rect 19901 21981 19935 22015
rect 22026 21981 22060 22015
rect 22293 21981 22327 22015
rect 3985 21913 4019 21947
rect 4185 21913 4219 21947
rect 2973 21845 3007 21879
rect 10333 21845 10367 21879
rect 17969 21845 18003 21879
rect 18797 21845 18831 21879
rect 20269 21845 20303 21879
rect 20453 21845 20487 21879
rect 20913 21845 20947 21879
rect 2145 21641 2179 21675
rect 2605 21641 2639 21675
rect 2973 21641 3007 21675
rect 4353 21641 4387 21675
rect 4905 21641 4939 21675
rect 5365 21641 5399 21675
rect 20821 21641 20855 21675
rect 1961 21573 1995 21607
rect 21097 21573 21131 21607
rect 21189 21573 21223 21607
rect 1593 21505 1627 21539
rect 2789 21505 2823 21539
rect 3065 21505 3099 21539
rect 4169 21505 4203 21539
rect 9965 21505 9999 21539
rect 10609 21505 10643 21539
rect 19901 21505 19935 21539
rect 21000 21505 21034 21539
rect 21317 21505 21351 21539
rect 21465 21505 21499 21539
rect 3525 21437 3559 21471
rect 19441 21437 19475 21471
rect 20361 21437 20395 21471
rect 20177 21369 20211 21403
rect 1961 21301 1995 21335
rect 10517 21301 10551 21335
rect 18705 21301 18739 21335
rect 22293 21301 22327 21335
rect 2145 21097 2179 21131
rect 2789 21097 2823 21131
rect 4077 21097 4111 21131
rect 4629 21097 4663 21131
rect 11713 21097 11747 21131
rect 20085 21097 20119 21131
rect 20269 21097 20303 21131
rect 22293 21097 22327 21131
rect 2605 21029 2639 21063
rect 1685 20961 1719 20995
rect 6653 20961 6687 20995
rect 10333 20961 10367 20995
rect 20913 20961 20947 20995
rect 1593 20893 1627 20927
rect 1869 20893 1903 20927
rect 1961 20893 1995 20927
rect 6745 20893 6779 20927
rect 10589 20893 10623 20927
rect 18889 20893 18923 20927
rect 19441 20893 19475 20927
rect 21169 20893 21203 20927
rect 2973 20825 3007 20859
rect 20237 20825 20271 20859
rect 20453 20825 20487 20859
rect 2773 20757 2807 20791
rect 7113 20757 7147 20791
rect 19625 20757 19659 20791
rect 1593 20553 1627 20587
rect 3249 20553 3283 20587
rect 14565 20553 14599 20587
rect 21297 20553 21331 20587
rect 21465 20553 21499 20587
rect 1777 20485 1811 20519
rect 7634 20485 7668 20519
rect 13860 20485 13894 20519
rect 21097 20485 21131 20519
rect 1961 20417 1995 20451
rect 3065 20417 3099 20451
rect 3709 20417 3743 20451
rect 7389 20417 7423 20451
rect 14933 20417 14967 20451
rect 19993 20417 20027 20451
rect 20637 20417 20671 20451
rect 14105 20349 14139 20383
rect 15025 20349 15059 20383
rect 12725 20281 12759 20315
rect 2421 20213 2455 20247
rect 8769 20213 8803 20247
rect 21281 20213 21315 20247
rect 22293 20213 22327 20247
rect 14289 20009 14323 20043
rect 21189 20009 21223 20043
rect 21925 20009 21959 20043
rect 22293 20009 22327 20043
rect 1593 19805 1627 19839
rect 2237 19805 2271 19839
rect 20729 19805 20763 19839
rect 21373 19805 21407 19839
rect 21833 19805 21867 19839
rect 2881 19737 2915 19771
rect 1777 19669 1811 19703
rect 2237 19465 2271 19499
rect 2421 19329 2455 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 12357 19329 12391 19363
rect 12516 19329 12550 19363
rect 13369 19329 13403 19363
rect 13553 19329 13587 19363
rect 21465 19329 21499 19363
rect 22293 19329 22327 19363
rect 12633 19261 12667 19295
rect 12909 19193 12943 19227
rect 22109 19193 22143 19227
rect 1593 19125 1627 19159
rect 2881 19125 2915 19159
rect 10977 19125 11011 19159
rect 1961 18921 1995 18955
rect 21557 18921 21591 18955
rect 2697 18853 2731 18887
rect 6929 18785 6963 18819
rect 2053 18717 2087 18751
rect 2513 18717 2547 18751
rect 3341 18717 3375 18751
rect 7021 18717 7055 18751
rect 22293 18717 22327 18751
rect 1593 18581 1627 18615
rect 3157 18581 3191 18615
rect 7389 18581 7423 18615
rect 2145 18377 2179 18411
rect 9229 18377 9263 18411
rect 1961 18309 1995 18343
rect 8094 18309 8128 18343
rect 2789 18241 2823 18275
rect 2973 18241 3007 18275
rect 3065 18241 3099 18275
rect 7849 18241 7883 18275
rect 1593 18173 1627 18207
rect 2605 18105 2639 18139
rect 22293 18105 22327 18139
rect 1961 18037 1995 18071
rect 3525 18037 3559 18071
rect 22109 17833 22143 17867
rect 1593 17629 1627 17663
rect 4169 17629 4203 17663
rect 4997 17629 5031 17663
rect 21649 17629 21683 17663
rect 22293 17629 22327 17663
rect 1838 17561 1872 17595
rect 3985 17561 4019 17595
rect 2973 17493 3007 17527
rect 4353 17493 4387 17527
rect 4813 17493 4847 17527
rect 2973 17289 3007 17323
rect 1860 17221 1894 17255
rect 3433 17153 3467 17187
rect 4537 17153 4571 17187
rect 4721 17153 4755 17187
rect 4813 17153 4847 17187
rect 1593 17085 1627 17119
rect 3709 17017 3743 17051
rect 5273 17017 5307 17051
rect 22293 17017 22327 17051
rect 3893 16949 3927 16983
rect 4353 16949 4387 16983
rect 4353 16745 4387 16779
rect 6009 16745 6043 16779
rect 4537 16677 4571 16711
rect 1593 16609 1627 16643
rect 3985 16609 4019 16643
rect 22293 16609 22327 16643
rect 1860 16541 1894 16575
rect 6653 16541 6687 16575
rect 6837 16541 6871 16575
rect 4997 16473 5031 16507
rect 5181 16473 5215 16507
rect 6193 16473 6227 16507
rect 2973 16405 3007 16439
rect 4353 16405 4387 16439
rect 5365 16405 5399 16439
rect 5825 16405 5859 16439
rect 5993 16405 6027 16439
rect 6653 16405 6687 16439
rect 1593 16201 1627 16235
rect 3433 16201 3467 16235
rect 22293 16201 22327 16235
rect 2728 16133 2762 16167
rect 6713 16133 6747 16167
rect 6929 16133 6963 16167
rect 2973 16065 3007 16099
rect 4557 16065 4591 16099
rect 21465 16065 21499 16099
rect 22109 16065 22143 16099
rect 4813 15997 4847 16031
rect 5733 15997 5767 16031
rect 5365 15929 5399 15963
rect 5273 15861 5307 15895
rect 6561 15861 6595 15895
rect 6745 15861 6779 15895
rect 4629 15657 4663 15691
rect 5089 15657 5123 15691
rect 5273 15657 5307 15691
rect 5917 15657 5951 15691
rect 6561 15657 6595 15691
rect 2605 15521 2639 15555
rect 1593 15453 1627 15487
rect 2421 15453 2455 15487
rect 2789 15453 2823 15487
rect 3065 15453 3099 15487
rect 3985 15453 4019 15487
rect 4078 15453 4112 15487
rect 4261 15453 4295 15487
rect 4491 15453 4525 15487
rect 6101 15453 6135 15487
rect 6745 15453 6779 15487
rect 7665 15453 7699 15487
rect 22293 15453 22327 15487
rect 4353 15385 4387 15419
rect 5257 15385 5291 15419
rect 5457 15385 5491 15419
rect 1869 15317 1903 15351
rect 7481 15317 7515 15351
rect 1593 15113 1627 15147
rect 3985 15113 4019 15147
rect 4905 15113 4939 15147
rect 5365 15113 5399 15147
rect 2728 15045 2762 15079
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 3709 14977 3743 15011
rect 3801 14977 3835 15011
rect 4445 14977 4479 15011
rect 5549 14977 5583 15011
rect 2973 14909 3007 14943
rect 4813 14841 4847 14875
rect 22293 14841 22327 14875
rect 4997 14569 5031 14603
rect 4813 14501 4847 14535
rect 2973 14433 3007 14467
rect 4353 14433 4387 14467
rect 2717 14365 2751 14399
rect 5641 14365 5675 14399
rect 3985 14297 4019 14331
rect 4169 14297 4203 14331
rect 5181 14297 5215 14331
rect 1593 14229 1627 14263
rect 4971 14229 5005 14263
rect 1961 14025 1995 14059
rect 2145 14025 2179 14059
rect 3157 14025 3191 14059
rect 3985 14025 4019 14059
rect 4537 14025 4571 14059
rect 2605 13889 2639 13923
rect 2881 13889 2915 13923
rect 2973 13889 3007 13923
rect 3617 13889 3651 13923
rect 3801 13889 3835 13923
rect 4445 13889 4479 13923
rect 2697 13821 2731 13855
rect 22293 13821 22327 13855
rect 1593 13753 1627 13787
rect 1961 13685 1995 13719
rect 1685 13481 1719 13515
rect 2145 13481 2179 13515
rect 2789 13481 2823 13515
rect 2973 13481 3007 13515
rect 4169 13481 4203 13515
rect 1593 13277 1627 13311
rect 1869 13277 1903 13311
rect 1961 13277 1995 13311
rect 3985 13277 4019 13311
rect 4629 13277 4663 13311
rect 22293 13277 22327 13311
rect 2631 13209 2665 13243
rect 2815 13141 2849 13175
rect 2605 12937 2639 12971
rect 1685 12801 1719 12835
rect 1777 12801 1811 12835
rect 2421 12801 2455 12835
rect 2605 12801 2639 12835
rect 3065 12801 3099 12835
rect 3893 12801 3927 12835
rect 4353 12801 4387 12835
rect 1961 12733 1995 12767
rect 3709 12597 3743 12631
rect 1777 12393 1811 12427
rect 2237 12393 2271 12427
rect 2973 12393 3007 12427
rect 1593 12189 1627 12223
rect 2881 12189 2915 12223
rect 22293 12189 22327 12223
rect 1685 11849 1719 11883
rect 1777 11713 1811 11747
rect 2237 11713 2271 11747
rect 22293 11577 22327 11611
rect 2881 11509 2915 11543
rect 1685 11305 1719 11339
rect 1593 11101 1627 11135
rect 1777 10761 1811 10795
rect 1593 10625 1627 10659
rect 2237 10625 2271 10659
rect 22293 10489 22327 10523
rect 1593 10013 1627 10047
rect 22293 10013 22327 10047
rect 1593 9333 1627 9367
rect 1593 9129 1627 9163
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 22293 8925 22327 8959
rect 22293 8313 22327 8347
rect 1593 7837 1627 7871
rect 22293 7225 22327 7259
rect 1593 7157 1627 7191
rect 22293 6749 22327 6783
rect 1869 6273 1903 6307
rect 1685 6069 1719 6103
rect 22293 5661 22327 5695
rect 1593 5117 1627 5151
rect 22293 5049 22327 5083
rect 22293 3961 22327 3995
rect 1593 3893 1627 3927
rect 1593 3485 1627 3519
rect 22293 3485 22327 3519
rect 1593 2805 1627 2839
rect 1593 2397 1627 2431
<< metal1 >>
rect 3970 27820 3976 27872
rect 4028 27860 4034 27872
rect 7466 27860 7472 27872
rect 4028 27832 7472 27860
rect 4028 27820 4034 27832
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 1104 27770 22816 27792
rect 1104 27718 3664 27770
rect 3716 27718 3728 27770
rect 3780 27718 3792 27770
rect 3844 27718 3856 27770
rect 3908 27718 3920 27770
rect 3972 27718 9092 27770
rect 9144 27718 9156 27770
rect 9208 27718 9220 27770
rect 9272 27718 9284 27770
rect 9336 27718 9348 27770
rect 9400 27718 14520 27770
rect 14572 27718 14584 27770
rect 14636 27718 14648 27770
rect 14700 27718 14712 27770
rect 14764 27718 14776 27770
rect 14828 27718 19948 27770
rect 20000 27718 20012 27770
rect 20064 27718 20076 27770
rect 20128 27718 20140 27770
rect 20192 27718 20204 27770
rect 20256 27718 22816 27770
rect 1104 27696 22816 27718
rect 4062 27616 4068 27668
rect 4120 27656 4126 27668
rect 7558 27656 7564 27668
rect 4120 27628 7564 27656
rect 4120 27616 4126 27628
rect 7558 27616 7564 27628
rect 7616 27616 7622 27668
rect 9309 27659 9367 27665
rect 9309 27625 9321 27659
rect 9355 27656 9367 27659
rect 11974 27656 11980 27668
rect 9355 27628 11980 27656
rect 9355 27625 9367 27628
rect 9309 27619 9367 27625
rect 11974 27616 11980 27628
rect 12032 27616 12038 27668
rect 12084 27628 12572 27656
rect 4709 27591 4767 27597
rect 4709 27557 4721 27591
rect 4755 27588 4767 27591
rect 6822 27588 6828 27600
rect 4755 27560 6828 27588
rect 4755 27557 4767 27560
rect 4709 27551 4767 27557
rect 6822 27548 6828 27560
rect 6880 27548 6886 27600
rect 8573 27591 8631 27597
rect 8573 27557 8585 27591
rect 8619 27588 8631 27591
rect 8619 27560 10180 27588
rect 8619 27557 8631 27560
rect 8573 27551 8631 27557
rect 3234 27520 3240 27532
rect 2746 27492 3240 27520
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27452 1639 27455
rect 1762 27452 1768 27464
rect 1627 27424 1768 27452
rect 1627 27421 1639 27424
rect 1581 27415 1639 27421
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 2225 27455 2283 27461
rect 2225 27421 2237 27455
rect 2271 27452 2283 27455
rect 2746 27452 2774 27492
rect 3234 27480 3240 27492
rect 3292 27480 3298 27532
rect 7193 27523 7251 27529
rect 7193 27520 7205 27523
rect 6472 27492 7205 27520
rect 2271 27424 2774 27452
rect 3053 27455 3111 27461
rect 2271 27421 2283 27424
rect 2225 27415 2283 27421
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 5169 27455 5227 27461
rect 5169 27421 5181 27455
rect 5215 27452 5227 27455
rect 5258 27452 5264 27464
rect 5215 27424 5264 27452
rect 5215 27421 5227 27424
rect 5169 27415 5227 27421
rect 3068 27384 3096 27415
rect 5258 27412 5264 27424
rect 5316 27412 5322 27464
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5718 27452 5724 27464
rect 5399 27424 5724 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 5813 27455 5871 27461
rect 5813 27421 5825 27455
rect 5859 27452 5871 27455
rect 6086 27452 6092 27464
rect 5859 27424 6092 27452
rect 5859 27421 5871 27424
rect 5813 27415 5871 27421
rect 6086 27412 6092 27424
rect 6144 27412 6150 27464
rect 6270 27384 6276 27396
rect 3068 27356 6276 27384
rect 6270 27344 6276 27356
rect 6328 27344 6334 27396
rect 1765 27319 1823 27325
rect 1765 27285 1777 27319
rect 1811 27316 1823 27319
rect 1854 27316 1860 27328
rect 1811 27288 1860 27316
rect 1811 27285 1823 27288
rect 1765 27279 1823 27285
rect 1854 27276 1860 27288
rect 1912 27276 1918 27328
rect 2406 27316 2412 27328
rect 2367 27288 2412 27316
rect 2406 27276 2412 27288
rect 2464 27276 2470 27328
rect 2958 27316 2964 27328
rect 2919 27288 2964 27316
rect 2958 27276 2964 27288
rect 3016 27276 3022 27328
rect 4062 27316 4068 27328
rect 4023 27288 4068 27316
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 5350 27316 5356 27328
rect 5311 27288 5356 27316
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 5997 27319 6055 27325
rect 5997 27285 6009 27319
rect 6043 27316 6055 27319
rect 6472 27316 6500 27492
rect 7193 27489 7205 27492
rect 7239 27489 7251 27523
rect 7193 27483 7251 27489
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 6730 27452 6736 27464
rect 6691 27424 6736 27452
rect 6549 27415 6607 27421
rect 6564 27384 6592 27415
rect 6730 27412 6736 27424
rect 6788 27412 6794 27464
rect 7208 27452 7236 27483
rect 10152 27452 10180 27560
rect 11072 27492 11744 27520
rect 11072 27452 11100 27492
rect 11716 27461 11744 27492
rect 7208 27424 10088 27452
rect 10152 27424 11100 27452
rect 11149 27455 11207 27461
rect 6822 27384 6828 27396
rect 6564 27356 6828 27384
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 6914 27344 6920 27396
rect 6972 27384 6978 27396
rect 7438 27387 7496 27393
rect 7438 27384 7450 27387
rect 6972 27356 7450 27384
rect 6972 27344 6978 27356
rect 7438 27353 7450 27356
rect 7484 27353 7496 27387
rect 10060 27384 10088 27424
rect 11149 27421 11161 27455
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 10318 27384 10324 27396
rect 10060 27356 10324 27384
rect 7438 27347 7496 27353
rect 10318 27344 10324 27356
rect 10376 27384 10382 27396
rect 10778 27384 10784 27396
rect 10376 27356 10784 27384
rect 10376 27344 10382 27356
rect 10778 27344 10784 27356
rect 10836 27344 10842 27396
rect 10882 27387 10940 27393
rect 10882 27353 10894 27387
rect 10928 27353 10940 27387
rect 10882 27347 10940 27353
rect 6043 27288 6500 27316
rect 6733 27319 6791 27325
rect 6043 27285 6055 27288
rect 5997 27279 6055 27285
rect 6733 27285 6745 27319
rect 6779 27316 6791 27319
rect 8386 27316 8392 27328
rect 6779 27288 8392 27316
rect 6779 27285 6791 27288
rect 6733 27279 6791 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 9769 27319 9827 27325
rect 9769 27285 9781 27319
rect 9815 27316 9827 27319
rect 10134 27316 10140 27328
rect 9815 27288 10140 27316
rect 9815 27285 9827 27288
rect 9769 27279 9827 27285
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 10686 27276 10692 27328
rect 10744 27316 10750 27328
rect 10897 27316 10925 27347
rect 11054 27344 11060 27396
rect 11112 27384 11118 27396
rect 11164 27384 11192 27415
rect 12084 27384 12112 27628
rect 12544 27588 12572 27628
rect 14458 27616 14464 27668
rect 14516 27656 14522 27668
rect 14516 27628 15516 27656
rect 14516 27616 14522 27628
rect 13998 27588 14004 27600
rect 12544 27560 14004 27588
rect 13998 27548 14004 27560
rect 14056 27548 14062 27600
rect 15488 27597 15516 27628
rect 15473 27591 15531 27597
rect 15473 27557 15485 27591
rect 15519 27557 15531 27591
rect 15473 27551 15531 27557
rect 16942 27548 16948 27600
rect 17000 27588 17006 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17000 27560 17509 27588
rect 17000 27548 17006 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 20073 27591 20131 27597
rect 20073 27588 20085 27591
rect 19484 27560 20085 27588
rect 19484 27548 19490 27560
rect 20073 27557 20085 27560
rect 20119 27557 20131 27591
rect 20073 27551 20131 27557
rect 20346 27548 20352 27600
rect 20404 27588 20410 27600
rect 20717 27591 20775 27597
rect 20717 27588 20729 27591
rect 20404 27560 20729 27588
rect 20404 27548 20410 27560
rect 20717 27557 20729 27560
rect 20763 27557 20775 27591
rect 20717 27551 20775 27557
rect 12710 27480 12716 27532
rect 12768 27520 12774 27532
rect 12768 27492 12813 27520
rect 12768 27480 12774 27492
rect 14182 27480 14188 27532
rect 14240 27520 14246 27532
rect 14240 27492 14596 27520
rect 14240 27480 14246 27492
rect 12526 27452 12532 27464
rect 12487 27424 12532 27452
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 12894 27452 12900 27464
rect 12855 27424 12900 27452
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 13078 27452 13084 27464
rect 13039 27424 13084 27452
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 13262 27412 13268 27464
rect 13320 27452 13326 27464
rect 14568 27461 14596 27492
rect 14642 27480 14648 27532
rect 14700 27520 14706 27532
rect 15381 27523 15439 27529
rect 14700 27492 14780 27520
rect 14700 27480 14706 27492
rect 14752 27461 14780 27492
rect 15381 27489 15393 27523
rect 15427 27489 15439 27523
rect 18785 27523 18843 27529
rect 18785 27520 18797 27523
rect 15381 27483 15439 27489
rect 18340 27492 18797 27520
rect 14456 27455 14514 27461
rect 14456 27452 14468 27455
rect 13320 27424 14468 27452
rect 13320 27412 13326 27424
rect 14456 27421 14468 27424
rect 14502 27421 14514 27455
rect 14456 27415 14514 27421
rect 14553 27455 14611 27461
rect 14553 27421 14565 27455
rect 14599 27421 14611 27455
rect 14752 27455 14831 27461
rect 14752 27424 14785 27455
rect 14553 27415 14611 27421
rect 14773 27421 14785 27424
rect 14819 27421 14831 27455
rect 14773 27415 14831 27421
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27452 14979 27455
rect 15396 27452 15424 27483
rect 17034 27452 17040 27464
rect 14967 27424 15424 27452
rect 16995 27424 17040 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18340 27461 18368 27492
rect 18785 27489 18797 27492
rect 18831 27489 18843 27523
rect 18785 27483 18843 27489
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 18012 27424 18337 27452
rect 18012 27412 18018 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18598 27412 18604 27464
rect 18656 27452 18662 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 18656 27424 19441 27452
rect 18656 27412 18662 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 20530 27412 20536 27464
rect 20588 27452 20594 27464
rect 21269 27455 21327 27461
rect 21269 27452 21281 27455
rect 20588 27424 21281 27452
rect 20588 27412 20594 27424
rect 21269 27421 21281 27424
rect 21315 27421 21327 27455
rect 22094 27452 22100 27464
rect 22055 27424 22100 27452
rect 21269 27415 21327 27421
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 11112 27356 12112 27384
rect 11112 27344 11118 27356
rect 13170 27344 13176 27396
rect 13228 27384 13234 27396
rect 14642 27384 14648 27396
rect 13228 27356 14504 27384
rect 14603 27356 14648 27384
rect 13228 27344 13234 27356
rect 10744 27288 10925 27316
rect 10744 27276 10750 27288
rect 11698 27276 11704 27328
rect 11756 27316 11762 27328
rect 11793 27319 11851 27325
rect 11793 27316 11805 27319
rect 11756 27288 11805 27316
rect 11756 27276 11762 27288
rect 11793 27285 11805 27288
rect 11839 27285 11851 27319
rect 11793 27279 11851 27285
rect 13446 27276 13452 27328
rect 13504 27316 13510 27328
rect 14277 27319 14335 27325
rect 14277 27316 14289 27319
rect 13504 27288 14289 27316
rect 13504 27276 13510 27288
rect 14277 27285 14289 27288
rect 14323 27285 14335 27319
rect 14476 27316 14504 27356
rect 14642 27344 14648 27356
rect 14700 27344 14706 27396
rect 15746 27344 15752 27396
rect 15804 27384 15810 27396
rect 15841 27387 15899 27393
rect 15841 27384 15853 27387
rect 15804 27356 15853 27384
rect 15804 27344 15810 27356
rect 15841 27353 15853 27356
rect 15887 27353 15899 27387
rect 15841 27347 15899 27353
rect 16853 27319 16911 27325
rect 16853 27316 16865 27319
rect 14476 27288 16865 27316
rect 14277 27279 14335 27285
rect 16853 27285 16865 27288
rect 16899 27285 16911 27319
rect 18138 27316 18144 27328
rect 18099 27288 18144 27316
rect 16853 27279 16911 27285
rect 18138 27276 18144 27288
rect 18196 27276 18202 27328
rect 21358 27316 21364 27328
rect 21319 27288 21364 27316
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 21818 27276 21824 27328
rect 21876 27316 21882 27328
rect 22189 27319 22247 27325
rect 22189 27316 22201 27319
rect 21876 27288 22201 27316
rect 21876 27276 21882 27288
rect 22189 27285 22201 27288
rect 22235 27285 22247 27319
rect 22189 27279 22247 27285
rect 1104 27226 22976 27248
rect 1104 27174 6378 27226
rect 6430 27174 6442 27226
rect 6494 27174 6506 27226
rect 6558 27174 6570 27226
rect 6622 27174 6634 27226
rect 6686 27174 11806 27226
rect 11858 27174 11870 27226
rect 11922 27174 11934 27226
rect 11986 27174 11998 27226
rect 12050 27174 12062 27226
rect 12114 27174 17234 27226
rect 17286 27174 17298 27226
rect 17350 27174 17362 27226
rect 17414 27174 17426 27226
rect 17478 27174 17490 27226
rect 17542 27174 22662 27226
rect 22714 27174 22726 27226
rect 22778 27174 22790 27226
rect 22842 27174 22854 27226
rect 22906 27174 22918 27226
rect 22970 27174 22976 27226
rect 1104 27152 22976 27174
rect 5350 27072 5356 27124
rect 5408 27112 5414 27124
rect 7167 27115 7225 27121
rect 7167 27112 7179 27115
rect 5408 27084 7179 27112
rect 5408 27072 5414 27084
rect 7167 27081 7179 27084
rect 7213 27081 7225 27115
rect 7929 27115 7987 27121
rect 7929 27112 7941 27115
rect 7167 27075 7225 27081
rect 7852 27084 7941 27112
rect 1578 27044 1584 27056
rect 1539 27016 1584 27044
rect 1578 27004 1584 27016
rect 1636 27004 1642 27056
rect 1797 27047 1855 27053
rect 1797 27013 1809 27047
rect 1843 27044 1855 27047
rect 3050 27044 3056 27056
rect 1843 27016 3056 27044
rect 1843 27013 1855 27016
rect 1797 27007 1855 27013
rect 3050 27004 3056 27016
rect 3108 27004 3114 27056
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 7006 27044 7012 27056
rect 4120 27016 7012 27044
rect 4120 27004 4126 27016
rect 2038 26936 2044 26988
rect 2096 26976 2102 26988
rect 2409 26979 2467 26985
rect 2409 26976 2421 26979
rect 2096 26948 2421 26976
rect 2096 26936 2102 26948
rect 2409 26945 2421 26948
rect 2455 26945 2467 26979
rect 2409 26939 2467 26945
rect 3510 26936 3516 26988
rect 3568 26976 3574 26988
rect 3789 26979 3847 26985
rect 3789 26976 3801 26979
rect 3568 26948 3801 26976
rect 3568 26936 3574 26948
rect 3789 26945 3801 26948
rect 3835 26945 3847 26979
rect 4522 26976 4528 26988
rect 4483 26948 4528 26976
rect 3789 26939 3847 26945
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 5166 26976 5172 26988
rect 5127 26948 5172 26976
rect 5166 26936 5172 26948
rect 5224 26936 5230 26988
rect 5828 26985 5856 27016
rect 7006 27004 7012 27016
rect 7064 27004 7070 27056
rect 7377 27047 7435 27053
rect 7377 27013 7389 27047
rect 7423 27044 7435 27047
rect 7650 27044 7656 27056
rect 7423 27016 7656 27044
rect 7423 27013 7435 27016
rect 7377 27007 7435 27013
rect 7650 27004 7656 27016
rect 7708 27004 7714 27056
rect 7742 27004 7748 27056
rect 7800 27044 7806 27056
rect 7852 27044 7880 27084
rect 7929 27081 7941 27084
rect 7975 27081 7987 27115
rect 7929 27075 7987 27081
rect 8018 27072 8024 27124
rect 8076 27112 8082 27124
rect 9950 27112 9956 27124
rect 8076 27084 9956 27112
rect 8076 27072 8082 27084
rect 9950 27072 9956 27084
rect 10008 27072 10014 27124
rect 10042 27072 10048 27124
rect 10100 27112 10106 27124
rect 11698 27112 11704 27124
rect 10100 27084 11704 27112
rect 10100 27072 10106 27084
rect 11698 27072 11704 27084
rect 11756 27072 11762 27124
rect 12526 27072 12532 27124
rect 12584 27112 12590 27124
rect 14093 27115 14151 27121
rect 14093 27112 14105 27115
rect 12584 27084 14105 27112
rect 12584 27072 12590 27084
rect 14093 27081 14105 27084
rect 14139 27081 14151 27115
rect 14550 27112 14556 27124
rect 14511 27084 14556 27112
rect 14093 27075 14151 27081
rect 14550 27072 14556 27084
rect 14608 27072 14614 27124
rect 20530 27112 20536 27124
rect 20491 27084 20536 27112
rect 20530 27072 20536 27084
rect 20588 27072 20594 27124
rect 7800 27016 7880 27044
rect 7800 27004 7806 27016
rect 8202 27004 8208 27056
rect 8260 27044 8266 27056
rect 9125 27047 9183 27053
rect 9125 27044 9137 27047
rect 8260 27016 9137 27044
rect 8260 27004 8266 27016
rect 9125 27013 9137 27016
rect 9171 27044 9183 27047
rect 10060 27044 10088 27072
rect 11974 27044 11980 27056
rect 9171 27016 10088 27044
rect 10704 27016 11980 27044
rect 9171 27013 9183 27016
rect 9125 27007 9183 27013
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 6822 26936 6828 26988
rect 6880 26976 6886 26988
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 6880 26948 7849 26976
rect 6880 26936 6886 26948
rect 7837 26945 7849 26948
rect 7883 26945 7895 26979
rect 7837 26939 7895 26945
rect 8113 26979 8171 26985
rect 8113 26945 8125 26979
rect 8159 26976 8171 26979
rect 10704 26976 10732 27016
rect 11974 27004 11980 27016
rect 12032 27004 12038 27056
rect 13078 27044 13084 27056
rect 12084 27016 13084 27044
rect 10870 26976 10876 26988
rect 10928 26985 10934 26988
rect 8159 26948 10732 26976
rect 10840 26948 10876 26976
rect 8159 26945 8171 26948
rect 8113 26939 8171 26945
rect 5258 26868 5264 26920
rect 5316 26908 5322 26920
rect 6638 26908 6644 26920
rect 5316 26880 6644 26908
rect 5316 26868 5322 26880
rect 6638 26868 6644 26880
rect 6696 26868 6702 26920
rect 7852 26908 7880 26939
rect 10870 26936 10876 26948
rect 10928 26939 10940 26985
rect 10928 26936 10934 26939
rect 11514 26936 11520 26988
rect 11572 26976 11578 26988
rect 12084 26976 12112 27016
rect 13078 27004 13084 27016
rect 13136 27044 13142 27056
rect 13136 27016 13584 27044
rect 13136 27004 13142 27016
rect 11572 26948 12112 26976
rect 12825 26979 12883 26985
rect 11572 26936 11578 26948
rect 12825 26945 12837 26979
rect 12871 26976 12883 26979
rect 13170 26976 13176 26988
rect 12871 26948 13176 26976
rect 12871 26945 12883 26948
rect 12825 26939 12883 26945
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 13556 26985 13584 27016
rect 13630 27004 13636 27056
rect 13688 27044 13694 27056
rect 15013 27047 15071 27053
rect 13688 27016 13952 27044
rect 13688 27004 13694 27016
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26945 13599 26979
rect 13814 26976 13820 26988
rect 13775 26948 13820 26976
rect 13541 26939 13599 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 13924 26985 13952 27016
rect 15013 27013 15025 27047
rect 15059 27044 15071 27047
rect 18138 27044 18144 27056
rect 15059 27016 18144 27044
rect 15059 27013 15071 27016
rect 15013 27007 15071 27013
rect 18138 27004 18144 27016
rect 18196 27004 18202 27056
rect 21910 27044 21916 27056
rect 19260 27016 21916 27044
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 15565 26979 15623 26985
rect 15565 26976 15577 26979
rect 14056 26948 15577 26976
rect 14056 26936 14062 26948
rect 15565 26945 15577 26948
rect 15611 26945 15623 26979
rect 15565 26939 15623 26945
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 19260 26985 19288 27016
rect 21910 27004 21916 27016
rect 21968 27004 21974 27056
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16632 26948 16865 26976
rect 16632 26936 16638 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 17773 26979 17831 26985
rect 17773 26945 17785 26979
rect 17819 26976 17831 26979
rect 19245 26979 19303 26985
rect 17819 26948 18184 26976
rect 17819 26945 17831 26948
rect 17773 26939 17831 26945
rect 18156 26920 18184 26948
rect 19245 26945 19257 26979
rect 19291 26945 19303 26979
rect 20346 26976 20352 26988
rect 20307 26948 20352 26976
rect 19245 26939 19303 26945
rect 20346 26936 20352 26948
rect 20404 26936 20410 26988
rect 22186 26976 22192 26988
rect 22147 26948 22192 26976
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 11149 26911 11207 26917
rect 7852 26880 9674 26908
rect 5997 26843 6055 26849
rect 5997 26809 6009 26843
rect 6043 26840 6055 26843
rect 8478 26840 8484 26852
rect 6043 26812 8484 26840
rect 6043 26809 6055 26812
rect 5997 26803 6055 26809
rect 8478 26800 8484 26812
rect 8536 26800 8542 26852
rect 8757 26843 8815 26849
rect 8757 26809 8769 26843
rect 8803 26840 8815 26843
rect 8938 26840 8944 26852
rect 8803 26812 8944 26840
rect 8803 26809 8815 26812
rect 8757 26803 8815 26809
rect 8938 26800 8944 26812
rect 8996 26800 9002 26852
rect 1670 26732 1676 26784
rect 1728 26772 1734 26784
rect 1765 26775 1823 26781
rect 1765 26772 1777 26775
rect 1728 26744 1777 26772
rect 1728 26732 1734 26744
rect 1765 26741 1777 26744
rect 1811 26741 1823 26775
rect 1765 26735 1823 26741
rect 1949 26775 2007 26781
rect 1949 26741 1961 26775
rect 1995 26772 2007 26775
rect 2498 26772 2504 26784
rect 1995 26744 2504 26772
rect 1995 26741 2007 26744
rect 1949 26735 2007 26741
rect 2498 26732 2504 26744
rect 2556 26732 2562 26784
rect 2593 26775 2651 26781
rect 2593 26741 2605 26775
rect 2639 26772 2651 26775
rect 2682 26772 2688 26784
rect 2639 26744 2688 26772
rect 2639 26741 2651 26744
rect 2593 26735 2651 26741
rect 2682 26732 2688 26744
rect 2740 26732 2746 26784
rect 2866 26732 2872 26784
rect 2924 26772 2930 26784
rect 3053 26775 3111 26781
rect 3053 26772 3065 26775
rect 2924 26744 3065 26772
rect 2924 26732 2930 26744
rect 3053 26741 3065 26744
rect 3099 26741 3111 26775
rect 5350 26772 5356 26784
rect 5311 26744 5356 26772
rect 3053 26735 3111 26741
rect 5350 26732 5356 26744
rect 5408 26732 5414 26784
rect 7006 26772 7012 26784
rect 6967 26744 7012 26772
rect 7006 26732 7012 26744
rect 7064 26732 7070 26784
rect 7193 26775 7251 26781
rect 7193 26741 7205 26775
rect 7239 26772 7251 26775
rect 7374 26772 7380 26784
rect 7239 26744 7380 26772
rect 7239 26741 7251 26744
rect 7193 26735 7251 26741
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 8297 26775 8355 26781
rect 8297 26741 8309 26775
rect 8343 26772 8355 26775
rect 9125 26775 9183 26781
rect 9125 26772 9137 26775
rect 8343 26744 9137 26772
rect 8343 26741 8355 26744
rect 8297 26735 8355 26741
rect 9125 26741 9137 26744
rect 9171 26741 9183 26775
rect 9125 26735 9183 26741
rect 9309 26775 9367 26781
rect 9309 26741 9321 26775
rect 9355 26772 9367 26775
rect 9490 26772 9496 26784
rect 9355 26744 9496 26772
rect 9355 26741 9367 26744
rect 9309 26735 9367 26741
rect 9490 26732 9496 26744
rect 9548 26732 9554 26784
rect 9646 26772 9674 26880
rect 11149 26877 11161 26911
rect 11195 26908 11207 26911
rect 11422 26908 11428 26920
rect 11195 26880 11428 26908
rect 11195 26877 11207 26880
rect 11149 26871 11207 26877
rect 11422 26868 11428 26880
rect 11480 26868 11486 26920
rect 13078 26868 13084 26920
rect 13136 26908 13142 26920
rect 13136 26880 15792 26908
rect 13136 26868 13142 26880
rect 14737 26843 14795 26849
rect 11164 26812 12204 26840
rect 9769 26775 9827 26781
rect 9769 26772 9781 26775
rect 9646 26744 9781 26772
rect 9769 26741 9781 26744
rect 9815 26772 9827 26775
rect 11164 26772 11192 26812
rect 9815 26744 11192 26772
rect 9815 26741 9827 26744
rect 9769 26735 9827 26741
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 11606 26772 11612 26784
rect 11296 26744 11612 26772
rect 11296 26732 11302 26744
rect 11606 26732 11612 26744
rect 11664 26772 11670 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 11664 26744 11713 26772
rect 11664 26732 11670 26744
rect 11701 26741 11713 26744
rect 11747 26741 11759 26775
rect 12176 26772 12204 26812
rect 14737 26809 14749 26843
rect 14783 26840 14795 26843
rect 14918 26840 14924 26852
rect 14783 26812 14924 26840
rect 14783 26809 14795 26812
rect 14737 26803 14795 26809
rect 14918 26800 14924 26812
rect 14976 26800 14982 26852
rect 15764 26849 15792 26880
rect 18138 26868 18144 26920
rect 18196 26868 18202 26920
rect 18601 26911 18659 26917
rect 18601 26877 18613 26911
rect 18647 26908 18659 26911
rect 20530 26908 20536 26920
rect 18647 26880 20536 26908
rect 18647 26877 18659 26880
rect 18601 26871 18659 26877
rect 20530 26868 20536 26880
rect 20588 26868 20594 26920
rect 15749 26843 15807 26849
rect 15749 26809 15761 26843
rect 15795 26840 15807 26843
rect 16209 26843 16267 26849
rect 16209 26840 16221 26843
rect 15795 26812 16221 26840
rect 15795 26809 15807 26812
rect 15749 26803 15807 26809
rect 16209 26809 16221 26812
rect 16255 26809 16267 26843
rect 16209 26803 16267 26809
rect 19889 26843 19947 26849
rect 19889 26809 19901 26843
rect 19935 26840 19947 26843
rect 21082 26840 21088 26852
rect 19935 26812 21088 26840
rect 19935 26809 19947 26812
rect 19889 26803 19947 26809
rect 21082 26800 21088 26812
rect 21140 26800 21146 26852
rect 12434 26772 12440 26784
rect 12176 26744 12440 26772
rect 11701 26735 11759 26741
rect 12434 26732 12440 26744
rect 12492 26732 12498 26784
rect 12894 26732 12900 26784
rect 12952 26772 12958 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 12952 26744 13645 26772
rect 12952 26732 12958 26744
rect 13633 26741 13645 26744
rect 13679 26741 13691 26775
rect 13633 26735 13691 26741
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 14642 26772 14648 26784
rect 13964 26744 14648 26772
rect 13964 26732 13970 26744
rect 14642 26732 14648 26744
rect 14700 26732 14706 26784
rect 17954 26772 17960 26784
rect 17915 26744 17960 26772
rect 17954 26732 17960 26744
rect 18012 26732 18018 26784
rect 21450 26772 21456 26784
rect 21411 26744 21456 26772
rect 21450 26732 21456 26744
rect 21508 26732 21514 26784
rect 21542 26732 21548 26784
rect 21600 26772 21606 26784
rect 22005 26775 22063 26781
rect 22005 26772 22017 26775
rect 21600 26744 22017 26772
rect 21600 26732 21606 26744
rect 22005 26741 22017 26744
rect 22051 26741 22063 26775
rect 22005 26735 22063 26741
rect 1104 26682 22816 26704
rect 1104 26630 3664 26682
rect 3716 26630 3728 26682
rect 3780 26630 3792 26682
rect 3844 26630 3856 26682
rect 3908 26630 3920 26682
rect 3972 26630 9092 26682
rect 9144 26630 9156 26682
rect 9208 26630 9220 26682
rect 9272 26630 9284 26682
rect 9336 26630 9348 26682
rect 9400 26630 14520 26682
rect 14572 26630 14584 26682
rect 14636 26630 14648 26682
rect 14700 26630 14712 26682
rect 14764 26630 14776 26682
rect 14828 26630 19948 26682
rect 20000 26630 20012 26682
rect 20064 26630 20076 26682
rect 20128 26630 20140 26682
rect 20192 26630 20204 26682
rect 20256 26630 22816 26682
rect 1104 26608 22816 26630
rect 2038 26568 2044 26580
rect 1999 26540 2044 26568
rect 2038 26528 2044 26540
rect 2096 26528 2102 26580
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 6730 26568 6736 26580
rect 4120 26540 6736 26568
rect 4120 26528 4126 26540
rect 6730 26528 6736 26540
rect 6788 26528 6794 26580
rect 6914 26568 6920 26580
rect 6875 26540 6920 26568
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 7374 26568 7380 26580
rect 7335 26540 7380 26568
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 7650 26528 7656 26580
rect 7708 26568 7714 26580
rect 8202 26568 8208 26580
rect 7708 26540 8208 26568
rect 7708 26528 7714 26540
rect 8202 26528 8208 26540
rect 8260 26528 8266 26580
rect 8389 26571 8447 26577
rect 8389 26537 8401 26571
rect 8435 26537 8447 26571
rect 8389 26531 8447 26537
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8619 26540 9996 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 1949 26503 2007 26509
rect 1949 26469 1961 26503
rect 1995 26500 2007 26503
rect 2222 26500 2228 26512
rect 1995 26472 2228 26500
rect 1995 26469 2007 26472
rect 1949 26463 2007 26469
rect 2222 26460 2228 26472
rect 2280 26460 2286 26512
rect 2774 26500 2780 26512
rect 2735 26472 2780 26500
rect 2774 26460 2780 26472
rect 2832 26460 2838 26512
rect 4617 26503 4675 26509
rect 4617 26469 4629 26503
rect 4663 26469 4675 26503
rect 4617 26463 4675 26469
rect 5629 26503 5687 26509
rect 5629 26469 5641 26503
rect 5675 26500 5687 26503
rect 7742 26500 7748 26512
rect 5675 26472 7748 26500
rect 5675 26469 5687 26472
rect 5629 26463 5687 26469
rect 2501 26435 2559 26441
rect 2501 26401 2513 26435
rect 2547 26432 2559 26435
rect 4632 26432 4660 26463
rect 7742 26460 7748 26472
rect 7800 26460 7806 26512
rect 8404 26500 8432 26531
rect 9674 26500 9680 26512
rect 8404 26472 9680 26500
rect 9674 26460 9680 26472
rect 9732 26460 9738 26512
rect 9766 26460 9772 26512
rect 9824 26460 9830 26512
rect 2547 26404 4660 26432
rect 6273 26435 6331 26441
rect 2547 26401 2559 26404
rect 2501 26395 2559 26401
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 8662 26432 8668 26444
rect 6319 26404 8668 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 8662 26392 8668 26404
rect 8720 26392 8726 26444
rect 9784 26432 9812 26460
rect 9140 26404 9812 26432
rect 9968 26432 9996 26540
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 10229 26571 10287 26577
rect 10100 26540 10145 26568
rect 10100 26528 10106 26540
rect 10229 26537 10241 26571
rect 10275 26568 10287 26571
rect 12802 26568 12808 26580
rect 10275 26540 12808 26568
rect 10275 26537 10287 26540
rect 10229 26531 10287 26537
rect 12802 26528 12808 26540
rect 12860 26528 12866 26580
rect 14458 26568 14464 26580
rect 14419 26540 14464 26568
rect 14458 26528 14464 26540
rect 14516 26528 14522 26580
rect 11974 26460 11980 26512
rect 12032 26500 12038 26512
rect 12069 26503 12127 26509
rect 12069 26500 12081 26503
rect 12032 26472 12081 26500
rect 12032 26460 12038 26472
rect 12069 26469 12081 26472
rect 12115 26469 12127 26503
rect 12069 26463 12127 26469
rect 12158 26460 12164 26512
rect 12216 26500 12222 26512
rect 12342 26500 12348 26512
rect 12216 26472 12348 26500
rect 12216 26460 12222 26472
rect 12342 26460 12348 26472
rect 12400 26500 12406 26512
rect 13078 26500 13084 26512
rect 12400 26472 13084 26500
rect 12400 26460 12406 26472
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 14274 26500 14280 26512
rect 14235 26472 14280 26500
rect 14274 26460 14280 26472
rect 14332 26460 14338 26512
rect 14366 26460 14372 26512
rect 14424 26500 14430 26512
rect 15105 26503 15163 26509
rect 15105 26500 15117 26503
rect 14424 26472 15117 26500
rect 14424 26460 14430 26472
rect 15105 26469 15117 26472
rect 15151 26469 15163 26503
rect 15105 26463 15163 26469
rect 9968 26404 10824 26432
rect 2406 26324 2412 26376
rect 2464 26364 2470 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 2464 26336 3985 26364
rect 2464 26324 2470 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4801 26367 4859 26373
rect 4801 26333 4813 26367
rect 4847 26333 4859 26367
rect 5442 26364 5448 26376
rect 5403 26336 5448 26364
rect 4801 26327 4859 26333
rect 1578 26296 1584 26308
rect 1539 26268 1584 26296
rect 1578 26256 1584 26268
rect 1636 26256 1642 26308
rect 2498 26256 2504 26308
rect 2556 26296 2562 26308
rect 3234 26296 3240 26308
rect 2556 26268 3240 26296
rect 2556 26256 2562 26268
rect 3234 26256 3240 26268
rect 3292 26256 3298 26308
rect 3326 26256 3332 26308
rect 3384 26296 3390 26308
rect 4065 26299 4123 26305
rect 4065 26296 4077 26299
rect 3384 26268 4077 26296
rect 3384 26256 3390 26268
rect 4065 26265 4077 26268
rect 4111 26265 4123 26299
rect 4065 26259 4123 26265
rect 4816 26240 4844 26327
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 5718 26324 5724 26376
rect 5776 26364 5782 26376
rect 6730 26364 6736 26376
rect 5776 26336 6592 26364
rect 6691 26336 6736 26364
rect 5776 26324 5782 26336
rect 2958 26228 2964 26240
rect 2919 26200 2964 26228
rect 2958 26188 2964 26200
rect 3016 26188 3022 26240
rect 3142 26188 3148 26240
rect 3200 26228 3206 26240
rect 4798 26228 4804 26240
rect 3200 26200 4804 26228
rect 3200 26188 3206 26200
rect 4798 26188 4804 26200
rect 4856 26188 4862 26240
rect 6564 26228 6592 26336
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 7745 26367 7803 26373
rect 7745 26364 7757 26367
rect 7484 26336 7757 26364
rect 6638 26256 6644 26308
rect 6696 26296 6702 26308
rect 7484 26296 7512 26336
rect 7745 26333 7757 26336
rect 7791 26364 7803 26367
rect 8846 26364 8852 26376
rect 7791 26336 8852 26364
rect 7791 26333 7803 26336
rect 7745 26327 7803 26333
rect 8846 26324 8852 26336
rect 8904 26324 8910 26376
rect 6696 26268 7512 26296
rect 7561 26299 7619 26305
rect 6696 26256 6702 26268
rect 7561 26265 7573 26299
rect 7607 26296 7619 26299
rect 8202 26296 8208 26308
rect 7607 26268 8064 26296
rect 8163 26268 8208 26296
rect 7607 26265 7619 26268
rect 7561 26259 7619 26265
rect 7576 26228 7604 26259
rect 6564 26200 7604 26228
rect 8036 26228 8064 26268
rect 8202 26256 8208 26268
rect 8260 26256 8266 26308
rect 8386 26256 8392 26308
rect 8444 26305 8450 26308
rect 8444 26299 8463 26305
rect 8451 26265 8463 26299
rect 9140 26296 9168 26404
rect 9677 26367 9735 26373
rect 9677 26333 9689 26367
rect 9723 26364 9735 26367
rect 9766 26364 9772 26376
rect 9723 26336 9772 26364
rect 9723 26333 9735 26336
rect 9677 26327 9735 26333
rect 9766 26324 9772 26336
rect 9824 26324 9830 26376
rect 10689 26367 10747 26373
rect 10689 26364 10701 26367
rect 10336 26336 10701 26364
rect 8444 26259 8463 26265
rect 8496 26268 9168 26296
rect 9217 26299 9275 26305
rect 8444 26256 8450 26259
rect 8496 26228 8524 26268
rect 9217 26265 9229 26299
rect 9263 26296 9275 26299
rect 10336 26296 10364 26336
rect 10689 26333 10701 26336
rect 10735 26333 10747 26367
rect 10796 26364 10824 26404
rect 11698 26392 11704 26444
rect 11756 26432 11762 26444
rect 13814 26432 13820 26444
rect 11756 26404 13820 26432
rect 11756 26392 11762 26404
rect 11238 26364 11244 26376
rect 10796 26336 11244 26364
rect 10689 26327 10747 26333
rect 9263 26268 10364 26296
rect 9263 26265 9275 26268
rect 9217 26259 9275 26265
rect 8036 26200 8524 26228
rect 9950 26188 9956 26240
rect 10008 26228 10014 26240
rect 10045 26231 10103 26237
rect 10045 26228 10057 26231
rect 10008 26200 10057 26228
rect 10008 26188 10014 26200
rect 10045 26197 10057 26200
rect 10091 26197 10103 26231
rect 10704 26228 10732 26327
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 12158 26364 12164 26376
rect 11480 26336 12164 26364
rect 11480 26324 11486 26336
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12820 26373 12848 26404
rect 13814 26392 13820 26404
rect 13872 26392 13878 26444
rect 17954 26392 17960 26444
rect 18012 26432 18018 26444
rect 21634 26432 21640 26444
rect 18012 26404 19564 26432
rect 21595 26404 21640 26432
rect 18012 26392 18018 26404
rect 12529 26367 12587 26373
rect 12529 26364 12541 26367
rect 12308 26336 12541 26364
rect 12308 26324 12314 26336
rect 12529 26333 12541 26336
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 12805 26367 12863 26373
rect 12805 26333 12817 26367
rect 12851 26333 12863 26367
rect 12805 26327 12863 26333
rect 12897 26367 12955 26373
rect 12897 26333 12909 26367
rect 12943 26333 12955 26367
rect 12897 26327 12955 26333
rect 10778 26256 10784 26308
rect 10836 26296 10842 26308
rect 10934 26299 10992 26305
rect 10934 26296 10946 26299
rect 10836 26268 10946 26296
rect 10836 26256 10842 26268
rect 10934 26265 10946 26268
rect 10980 26265 10992 26299
rect 11440 26296 11468 26324
rect 12710 26296 12716 26308
rect 10934 26259 10992 26265
rect 11072 26268 11468 26296
rect 12671 26268 12716 26296
rect 11072 26228 11100 26268
rect 12710 26256 12716 26268
rect 12768 26256 12774 26308
rect 12912 26296 12940 26327
rect 12986 26324 12992 26376
rect 13044 26364 13050 26376
rect 13538 26364 13544 26376
rect 13044 26336 13544 26364
rect 13044 26324 13050 26336
rect 13538 26324 13544 26336
rect 13596 26364 13602 26376
rect 13725 26367 13783 26373
rect 13725 26364 13737 26367
rect 13596 26336 13737 26364
rect 13596 26324 13602 26336
rect 13725 26333 13737 26336
rect 13771 26333 13783 26367
rect 13725 26327 13783 26333
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 15933 26367 15991 26373
rect 15933 26364 15945 26367
rect 15344 26336 15945 26364
rect 15344 26324 15350 26336
rect 15933 26333 15945 26336
rect 15979 26364 15991 26367
rect 16393 26367 16451 26373
rect 16393 26364 16405 26367
rect 15979 26336 16405 26364
rect 15979 26333 15991 26336
rect 15933 26327 15991 26333
rect 16393 26333 16405 26336
rect 16439 26333 16451 26367
rect 16393 26327 16451 26333
rect 18877 26367 18935 26373
rect 18877 26333 18889 26367
rect 18923 26364 18935 26367
rect 19426 26364 19432 26376
rect 18923 26336 19432 26364
rect 18923 26333 18935 26336
rect 18877 26327 18935 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19536 26373 19564 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 20349 26367 20407 26373
rect 20349 26333 20361 26367
rect 20395 26364 20407 26367
rect 20622 26364 20628 26376
rect 20395 26336 20628 26364
rect 20395 26333 20407 26336
rect 20349 26327 20407 26333
rect 20622 26324 20628 26336
rect 20680 26324 20686 26376
rect 13170 26296 13176 26308
rect 12912 26268 13176 26296
rect 13170 26256 13176 26268
rect 13228 26296 13234 26308
rect 13630 26296 13636 26308
rect 13228 26268 13636 26296
rect 13228 26256 13234 26268
rect 13630 26256 13636 26268
rect 13688 26256 13694 26308
rect 14182 26256 14188 26308
rect 14240 26296 14246 26308
rect 14429 26299 14487 26305
rect 14429 26296 14441 26299
rect 14240 26268 14441 26296
rect 14240 26256 14246 26268
rect 14429 26265 14441 26268
rect 14475 26265 14487 26299
rect 14429 26259 14487 26265
rect 14645 26299 14703 26305
rect 14645 26265 14657 26299
rect 14691 26296 14703 26299
rect 14918 26296 14924 26308
rect 14691 26268 14924 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 10704 26200 11100 26228
rect 10045 26191 10103 26197
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 13081 26231 13139 26237
rect 13081 26228 13093 26231
rect 12584 26200 13093 26228
rect 12584 26188 12590 26200
rect 13081 26197 13093 26200
rect 13127 26197 13139 26231
rect 13081 26191 13139 26197
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 13541 26231 13599 26237
rect 13541 26228 13553 26231
rect 13412 26200 13553 26228
rect 13412 26188 13418 26200
rect 13541 26197 13553 26200
rect 13587 26197 13599 26231
rect 13541 26191 13599 26197
rect 14274 26188 14280 26240
rect 14332 26228 14338 26240
rect 14660 26228 14688 26259
rect 14918 26256 14924 26268
rect 14976 26256 14982 26308
rect 18138 26296 18144 26308
rect 18099 26268 18144 26296
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 19613 26299 19671 26305
rect 19613 26296 19625 26299
rect 19536 26268 19625 26296
rect 19536 26240 19564 26268
rect 19613 26265 19625 26268
rect 19659 26265 19671 26299
rect 20806 26296 20812 26308
rect 20767 26268 20812 26296
rect 19613 26259 19671 26265
rect 20806 26256 20812 26268
rect 20864 26256 20870 26308
rect 20898 26256 20904 26308
rect 20956 26296 20962 26308
rect 20993 26299 21051 26305
rect 20993 26296 21005 26299
rect 20956 26268 21005 26296
rect 20956 26256 20962 26268
rect 20993 26265 21005 26268
rect 21039 26265 21051 26299
rect 20993 26259 21051 26265
rect 21177 26299 21235 26305
rect 21177 26265 21189 26299
rect 21223 26296 21235 26299
rect 21266 26296 21272 26308
rect 21223 26268 21272 26296
rect 21223 26265 21235 26268
rect 21177 26259 21235 26265
rect 21266 26256 21272 26268
rect 21324 26256 21330 26308
rect 21634 26256 21640 26308
rect 21692 26296 21698 26308
rect 21821 26299 21879 26305
rect 21821 26296 21833 26299
rect 21692 26268 21833 26296
rect 21692 26256 21698 26268
rect 21821 26265 21833 26268
rect 21867 26265 21879 26299
rect 21821 26259 21879 26265
rect 21910 26256 21916 26308
rect 21968 26296 21974 26308
rect 22005 26299 22063 26305
rect 22005 26296 22017 26299
rect 21968 26268 22017 26296
rect 21968 26256 21974 26268
rect 22005 26265 22017 26268
rect 22051 26265 22063 26299
rect 22005 26259 22063 26265
rect 15746 26228 15752 26240
rect 14332 26200 14688 26228
rect 15707 26200 15752 26228
rect 14332 26188 14338 26200
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 19518 26188 19524 26240
rect 19576 26188 19582 26240
rect 1104 26138 22976 26160
rect 1104 26086 6378 26138
rect 6430 26086 6442 26138
rect 6494 26086 6506 26138
rect 6558 26086 6570 26138
rect 6622 26086 6634 26138
rect 6686 26086 11806 26138
rect 11858 26086 11870 26138
rect 11922 26086 11934 26138
rect 11986 26086 11998 26138
rect 12050 26086 12062 26138
rect 12114 26086 17234 26138
rect 17286 26086 17298 26138
rect 17350 26086 17362 26138
rect 17414 26086 17426 26138
rect 17478 26086 17490 26138
rect 17542 26086 22662 26138
rect 22714 26086 22726 26138
rect 22778 26086 22790 26138
rect 22842 26086 22854 26138
rect 22906 26086 22918 26138
rect 22970 26086 22976 26138
rect 1104 26064 22976 26086
rect 1578 25984 1584 26036
rect 1636 26024 1642 26036
rect 2685 26027 2743 26033
rect 2685 26024 2697 26027
rect 1636 25996 2697 26024
rect 1636 25984 1642 25996
rect 2685 25993 2697 25996
rect 2731 25993 2743 26027
rect 2685 25987 2743 25993
rect 1949 25959 2007 25965
rect 1949 25925 1961 25959
rect 1995 25956 2007 25959
rect 2222 25956 2228 25968
rect 1995 25928 2228 25956
rect 1995 25925 2007 25928
rect 1949 25919 2007 25925
rect 2222 25916 2228 25928
rect 2280 25916 2286 25968
rect 2700 25956 2728 25987
rect 3234 25984 3240 26036
rect 3292 26024 3298 26036
rect 5534 26024 5540 26036
rect 3292 25996 5540 26024
rect 3292 25984 3298 25996
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 10134 26024 10140 26036
rect 9646 25996 10140 26024
rect 2774 25956 2780 25968
rect 2700 25928 2780 25956
rect 2774 25916 2780 25928
rect 2832 25956 2838 25968
rect 9122 25965 9128 25968
rect 3697 25959 3755 25965
rect 3697 25956 3709 25959
rect 2832 25928 3709 25956
rect 2832 25916 2838 25928
rect 3697 25925 3709 25928
rect 3743 25956 3755 25959
rect 9109 25959 9128 25965
rect 9109 25956 9121 25959
rect 3743 25928 4384 25956
rect 3743 25925 3755 25928
rect 3697 25919 3755 25925
rect 1670 25848 1676 25900
rect 1728 25888 1734 25900
rect 2406 25888 2412 25900
rect 1728 25860 2412 25888
rect 1728 25848 1734 25860
rect 2406 25848 2412 25860
rect 2464 25888 2470 25900
rect 2593 25891 2651 25897
rect 2593 25888 2605 25891
rect 2464 25860 2605 25888
rect 2464 25848 2470 25860
rect 2593 25857 2605 25860
rect 2639 25857 2651 25891
rect 2593 25851 2651 25857
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25888 2927 25891
rect 3050 25888 3056 25900
rect 2915 25860 3056 25888
rect 2915 25857 2927 25860
rect 2869 25851 2927 25857
rect 2608 25820 2636 25851
rect 3050 25848 3056 25860
rect 3108 25848 3114 25900
rect 3881 25891 3939 25897
rect 3881 25857 3893 25891
rect 3927 25888 3939 25891
rect 4246 25888 4252 25900
rect 3927 25860 4252 25888
rect 3927 25857 3939 25860
rect 3881 25851 3939 25857
rect 3896 25820 3924 25851
rect 4246 25848 4252 25860
rect 4304 25848 4310 25900
rect 4356 25897 4384 25928
rect 8312 25928 9121 25956
rect 4341 25891 4399 25897
rect 4341 25857 4353 25891
rect 4387 25857 4399 25891
rect 4341 25851 4399 25857
rect 4430 25848 4436 25900
rect 4488 25888 4494 25900
rect 4525 25891 4583 25897
rect 4525 25888 4537 25891
rect 4488 25860 4537 25888
rect 4488 25848 4494 25860
rect 4525 25857 4537 25860
rect 4571 25857 4583 25891
rect 4525 25851 4583 25857
rect 6178 25848 6184 25900
rect 6236 25888 6242 25900
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 6236 25860 6561 25888
rect 6236 25848 6242 25860
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 7006 25848 7012 25900
rect 7064 25888 7070 25900
rect 8312 25897 8340 25928
rect 9109 25925 9121 25928
rect 9109 25919 9128 25925
rect 9122 25916 9128 25919
rect 9180 25916 9186 25968
rect 9309 25959 9367 25965
rect 9309 25925 9321 25959
rect 9355 25956 9367 25959
rect 9646 25956 9674 25996
rect 10134 25984 10140 25996
rect 10192 26024 10198 26036
rect 10192 25996 10977 26024
rect 10192 25984 10198 25996
rect 10949 25956 10977 25996
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 11149 26027 11207 26033
rect 11149 26024 11161 26027
rect 11112 25996 11161 26024
rect 11112 25984 11118 25996
rect 11149 25993 11161 25996
rect 11195 26024 11207 26027
rect 11698 26024 11704 26036
rect 11195 25996 11704 26024
rect 11195 25993 11207 25996
rect 11149 25987 11207 25993
rect 11698 25984 11704 25996
rect 11756 25984 11762 26036
rect 12250 26024 12256 26036
rect 11900 25996 12256 26024
rect 11422 25956 11428 25968
rect 9355 25928 9674 25956
rect 9784 25928 10180 25956
rect 10949 25928 11428 25956
rect 9355 25925 9367 25928
rect 9309 25919 9367 25925
rect 7469 25891 7527 25897
rect 7469 25888 7481 25891
rect 7064 25860 7481 25888
rect 7064 25848 7070 25860
rect 7469 25857 7481 25860
rect 7515 25857 7527 25891
rect 7469 25851 7527 25857
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 8297 25851 8355 25857
rect 2608 25792 3924 25820
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 5629 25823 5687 25829
rect 5629 25820 5641 25823
rect 4120 25792 5641 25820
rect 4120 25780 4126 25792
rect 5629 25789 5641 25792
rect 5675 25789 5687 25823
rect 5629 25783 5687 25789
rect 8113 25823 8171 25829
rect 8113 25789 8125 25823
rect 8159 25820 8171 25823
rect 9324 25820 9352 25919
rect 9784 25897 9812 25928
rect 9776 25891 9834 25897
rect 9776 25857 9788 25891
rect 9822 25857 9834 25891
rect 10025 25891 10083 25897
rect 10025 25888 10037 25891
rect 9968 25886 10037 25888
rect 9776 25851 9834 25857
rect 9876 25860 10037 25886
rect 9876 25858 9996 25860
rect 8159 25792 9352 25820
rect 8159 25789 8171 25792
rect 8113 25783 8171 25789
rect 9674 25780 9680 25832
rect 9732 25820 9738 25832
rect 9876 25820 9904 25858
rect 10025 25857 10037 25860
rect 10071 25857 10083 25891
rect 10152 25888 10180 25928
rect 11422 25916 11428 25928
rect 11480 25956 11486 25968
rect 11900 25956 11928 25996
rect 12250 25984 12256 25996
rect 12308 25984 12314 26036
rect 13173 26027 13231 26033
rect 13173 25993 13185 26027
rect 13219 26024 13231 26027
rect 13906 26024 13912 26036
rect 13219 25996 13912 26024
rect 13219 25993 13231 25996
rect 13173 25987 13231 25993
rect 13906 25984 13912 25996
rect 13964 25984 13970 26036
rect 18138 25984 18144 26036
rect 18196 26024 18202 26036
rect 22462 26024 22468 26036
rect 18196 25996 22468 26024
rect 18196 25984 18202 25996
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 12158 25956 12164 25968
rect 11480 25928 11928 25956
rect 11992 25928 12164 25956
rect 11480 25916 11486 25928
rect 10318 25888 10324 25900
rect 10152 25860 10324 25888
rect 10025 25851 10083 25857
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 10502 25848 10508 25900
rect 10560 25888 10566 25900
rect 11716 25897 11744 25928
rect 11992 25897 12020 25928
rect 12158 25916 12164 25928
rect 12216 25916 12222 25968
rect 15746 25956 15752 25968
rect 12728 25928 15752 25956
rect 12728 25897 12756 25928
rect 15746 25916 15752 25928
rect 15804 25916 15810 25968
rect 11701 25891 11759 25897
rect 10560 25860 10824 25888
rect 10560 25848 10566 25860
rect 9732 25792 9904 25820
rect 9732 25780 9738 25792
rect 1581 25755 1639 25761
rect 1581 25721 1593 25755
rect 1627 25752 1639 25755
rect 2038 25752 2044 25764
rect 1627 25724 2044 25752
rect 1627 25721 1639 25724
rect 1581 25715 1639 25721
rect 2038 25712 2044 25724
rect 2096 25712 2102 25764
rect 2130 25712 2136 25764
rect 2188 25752 2194 25764
rect 2188 25724 2233 25752
rect 2188 25712 2194 25724
rect 3418 25712 3424 25764
rect 3476 25752 3482 25764
rect 4985 25755 5043 25761
rect 4985 25752 4997 25755
rect 3476 25724 4997 25752
rect 3476 25712 3482 25724
rect 4985 25721 4997 25724
rect 5031 25721 5043 25755
rect 4985 25715 5043 25721
rect 8846 25712 8852 25764
rect 8904 25752 8910 25764
rect 8941 25755 8999 25761
rect 8941 25752 8953 25755
rect 8904 25724 8953 25752
rect 8904 25712 8910 25724
rect 8941 25721 8953 25724
rect 8987 25721 8999 25755
rect 9766 25752 9772 25764
rect 8941 25715 8999 25721
rect 9048 25724 9772 25752
rect 1946 25684 1952 25696
rect 1907 25656 1952 25684
rect 1946 25644 1952 25656
rect 2004 25644 2010 25696
rect 3050 25684 3056 25696
rect 3011 25656 3056 25684
rect 3050 25644 3056 25656
rect 3108 25644 3114 25696
rect 3234 25644 3240 25696
rect 3292 25684 3298 25696
rect 3513 25687 3571 25693
rect 3513 25684 3525 25687
rect 3292 25656 3525 25684
rect 3292 25644 3298 25656
rect 3513 25653 3525 25656
rect 3559 25653 3571 25687
rect 3513 25647 3571 25653
rect 3602 25644 3608 25696
rect 3660 25684 3666 25696
rect 4433 25687 4491 25693
rect 4433 25684 4445 25687
rect 3660 25656 4445 25684
rect 3660 25644 3666 25656
rect 4433 25653 4445 25656
rect 4479 25653 4491 25687
rect 7650 25684 7656 25696
rect 7611 25656 7656 25684
rect 4433 25647 4491 25653
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 8481 25687 8539 25693
rect 8481 25653 8493 25687
rect 8527 25684 8539 25687
rect 9048 25684 9076 25724
rect 9766 25712 9772 25724
rect 9824 25712 9830 25764
rect 10796 25752 10824 25860
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25857 12035 25891
rect 11977 25851 12035 25857
rect 12069 25891 12127 25897
rect 12069 25857 12081 25891
rect 12115 25888 12127 25891
rect 12713 25891 12771 25897
rect 12115 25860 12434 25888
rect 12115 25857 12127 25860
rect 12069 25851 12127 25857
rect 12406 25820 12434 25860
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 13262 25888 13268 25900
rect 12713 25851 12771 25857
rect 13096 25860 13268 25888
rect 13096 25820 13124 25860
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13817 25891 13875 25897
rect 13817 25857 13829 25891
rect 13863 25857 13875 25891
rect 13817 25851 13875 25857
rect 14001 25891 14059 25897
rect 14001 25857 14013 25891
rect 14047 25888 14059 25891
rect 14366 25888 14372 25900
rect 14047 25860 14372 25888
rect 14047 25857 14059 25860
rect 14001 25851 14059 25857
rect 12406 25792 13124 25820
rect 13280 25792 13676 25820
rect 13280 25752 13308 25792
rect 13648 25761 13676 25792
rect 10796 25724 13308 25752
rect 13633 25755 13691 25761
rect 13633 25721 13645 25755
rect 13679 25721 13691 25755
rect 13832 25752 13860 25851
rect 14366 25848 14372 25860
rect 14424 25848 14430 25900
rect 18693 25891 18751 25897
rect 18693 25857 18705 25891
rect 18739 25888 18751 25891
rect 19153 25891 19211 25897
rect 19153 25888 19165 25891
rect 18739 25860 19165 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 19153 25857 19165 25860
rect 19199 25888 19211 25891
rect 19426 25888 19432 25900
rect 19199 25860 19432 25888
rect 19199 25857 19211 25860
rect 19153 25851 19211 25857
rect 19426 25848 19432 25860
rect 19484 25848 19490 25900
rect 19702 25848 19708 25900
rect 19760 25888 19766 25900
rect 19797 25891 19855 25897
rect 19797 25888 19809 25891
rect 19760 25860 19809 25888
rect 19760 25848 19766 25860
rect 19797 25857 19809 25860
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 20346 25848 20352 25900
rect 20404 25888 20410 25900
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20404 25860 20453 25888
rect 20404 25848 20410 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 20441 25851 20499 25857
rect 20548 25860 21281 25888
rect 13906 25780 13912 25832
rect 13964 25820 13970 25832
rect 14461 25823 14519 25829
rect 14461 25820 14473 25823
rect 13964 25792 14473 25820
rect 13964 25780 13970 25792
rect 14461 25789 14473 25792
rect 14507 25789 14519 25823
rect 14461 25783 14519 25789
rect 19886 25780 19892 25832
rect 19944 25820 19950 25832
rect 20548 25820 20576 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 21726 25848 21732 25900
rect 21784 25888 21790 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21784 25860 22017 25888
rect 21784 25848 21790 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 21082 25820 21088 25832
rect 19944 25792 20576 25820
rect 21043 25792 21088 25820
rect 19944 25780 19950 25792
rect 21082 25780 21088 25792
rect 21140 25780 21146 25832
rect 14274 25752 14280 25764
rect 13832 25724 14280 25752
rect 13633 25715 13691 25721
rect 14274 25712 14280 25724
rect 14332 25712 14338 25764
rect 19337 25755 19395 25761
rect 19337 25721 19349 25755
rect 19383 25752 19395 25755
rect 22094 25752 22100 25764
rect 19383 25724 22100 25752
rect 19383 25721 19395 25724
rect 19337 25715 19395 25721
rect 22094 25712 22100 25724
rect 22152 25712 22158 25764
rect 8527 25656 9076 25684
rect 9125 25687 9183 25693
rect 8527 25653 8539 25656
rect 8481 25647 8539 25653
rect 9125 25653 9137 25687
rect 9171 25684 9183 25687
rect 11054 25684 11060 25696
rect 9171 25656 11060 25684
rect 9171 25653 9183 25656
rect 9125 25647 9183 25653
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 11790 25684 11796 25696
rect 11751 25656 11796 25684
rect 11790 25644 11796 25656
rect 11848 25644 11854 25696
rect 12250 25684 12256 25696
rect 12211 25656 12256 25684
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 12434 25644 12440 25696
rect 12492 25684 12498 25696
rect 12989 25687 13047 25693
rect 12989 25684 13001 25687
rect 12492 25656 13001 25684
rect 12492 25644 12498 25656
rect 12989 25653 13001 25656
rect 13035 25684 13047 25687
rect 13078 25684 13084 25696
rect 13035 25656 13084 25684
rect 13035 25653 13047 25656
rect 12989 25647 13047 25653
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 13538 25644 13544 25696
rect 13596 25684 13602 25696
rect 15197 25687 15255 25693
rect 15197 25684 15209 25687
rect 13596 25656 15209 25684
rect 13596 25644 13602 25656
rect 15197 25653 15209 25656
rect 15243 25653 15255 25687
rect 15197 25647 15255 25653
rect 19981 25687 20039 25693
rect 19981 25653 19993 25687
rect 20027 25684 20039 25687
rect 20530 25684 20536 25696
rect 20027 25656 20536 25684
rect 20027 25653 20039 25656
rect 19981 25647 20039 25653
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 20625 25687 20683 25693
rect 20625 25653 20637 25687
rect 20671 25684 20683 25687
rect 21174 25684 21180 25696
rect 20671 25656 21180 25684
rect 20671 25653 20683 25656
rect 20625 25647 20683 25653
rect 21174 25644 21180 25656
rect 21232 25644 21238 25696
rect 21266 25644 21272 25696
rect 21324 25684 21330 25696
rect 21453 25687 21511 25693
rect 21453 25684 21465 25687
rect 21324 25656 21465 25684
rect 21324 25644 21330 25656
rect 21453 25653 21465 25656
rect 21499 25653 21511 25687
rect 21453 25647 21511 25653
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 22189 25687 22247 25693
rect 22189 25684 22201 25687
rect 22060 25656 22201 25684
rect 22060 25644 22066 25656
rect 22189 25653 22201 25656
rect 22235 25653 22247 25687
rect 22189 25647 22247 25653
rect 1104 25594 22816 25616
rect 1104 25542 3664 25594
rect 3716 25542 3728 25594
rect 3780 25542 3792 25594
rect 3844 25542 3856 25594
rect 3908 25542 3920 25594
rect 3972 25542 9092 25594
rect 9144 25542 9156 25594
rect 9208 25542 9220 25594
rect 9272 25542 9284 25594
rect 9336 25542 9348 25594
rect 9400 25542 14520 25594
rect 14572 25542 14584 25594
rect 14636 25542 14648 25594
rect 14700 25542 14712 25594
rect 14764 25542 14776 25594
rect 14828 25542 19948 25594
rect 20000 25542 20012 25594
rect 20064 25542 20076 25594
rect 20128 25542 20140 25594
rect 20192 25542 20204 25594
rect 20256 25542 22816 25594
rect 1104 25520 22816 25542
rect 1578 25480 1584 25492
rect 1539 25452 1584 25480
rect 1578 25440 1584 25452
rect 1636 25440 1642 25492
rect 2314 25440 2320 25492
rect 2372 25480 2378 25492
rect 6181 25483 6239 25489
rect 6181 25480 6193 25483
rect 2372 25452 6193 25480
rect 2372 25440 2378 25452
rect 6181 25449 6193 25452
rect 6227 25449 6239 25483
rect 6181 25443 6239 25449
rect 6270 25440 6276 25492
rect 6328 25480 6334 25492
rect 6825 25483 6883 25489
rect 6825 25480 6837 25483
rect 6328 25452 6837 25480
rect 6328 25440 6334 25452
rect 6825 25449 6837 25452
rect 6871 25449 6883 25483
rect 7834 25480 7840 25492
rect 7795 25452 7840 25480
rect 6825 25443 6883 25449
rect 7834 25440 7840 25452
rect 7892 25440 7898 25492
rect 8481 25483 8539 25489
rect 8481 25449 8493 25483
rect 8527 25480 8539 25483
rect 11790 25480 11796 25492
rect 8527 25452 11796 25480
rect 8527 25449 8539 25452
rect 8481 25443 8539 25449
rect 11790 25440 11796 25452
rect 11848 25480 11854 25492
rect 13262 25480 13268 25492
rect 11848 25452 12434 25480
rect 13223 25452 13268 25480
rect 11848 25440 11854 25452
rect 4246 25412 4252 25424
rect 4207 25384 4252 25412
rect 4246 25372 4252 25384
rect 4304 25412 4310 25424
rect 4522 25412 4528 25424
rect 4304 25384 4528 25412
rect 4304 25372 4310 25384
rect 4522 25372 4528 25384
rect 4580 25372 4586 25424
rect 7650 25372 7656 25424
rect 7708 25412 7714 25424
rect 12406 25412 12434 25452
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 19334 25440 19340 25492
rect 19392 25480 19398 25492
rect 19794 25480 19800 25492
rect 19392 25452 19800 25480
rect 19392 25440 19398 25452
rect 19794 25440 19800 25452
rect 19852 25480 19858 25492
rect 20073 25483 20131 25489
rect 20073 25480 20085 25483
rect 19852 25452 20085 25480
rect 19852 25440 19858 25452
rect 20073 25449 20085 25452
rect 20119 25449 20131 25483
rect 20073 25443 20131 25449
rect 20257 25483 20315 25489
rect 20257 25449 20269 25483
rect 20303 25449 20315 25483
rect 20257 25443 20315 25449
rect 12710 25412 12716 25424
rect 7708 25384 10456 25412
rect 12406 25384 12716 25412
rect 7708 25372 7714 25384
rect 5537 25347 5595 25353
rect 5537 25344 5549 25347
rect 4264 25316 5549 25344
rect 4264 25288 4292 25316
rect 5537 25313 5549 25316
rect 5583 25313 5595 25347
rect 5537 25307 5595 25313
rect 9766 25304 9772 25356
rect 9824 25304 9830 25356
rect 10428 25344 10456 25384
rect 12710 25372 12716 25384
rect 12768 25372 12774 25424
rect 20272 25412 20300 25443
rect 20438 25440 20444 25492
rect 20496 25480 20502 25492
rect 20898 25480 20904 25492
rect 20496 25452 20904 25480
rect 20496 25440 20502 25452
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 20714 25412 20720 25424
rect 20272 25384 20720 25412
rect 20714 25372 20720 25384
rect 20772 25372 20778 25424
rect 10428 25316 10548 25344
rect 2682 25276 2688 25288
rect 2740 25285 2746 25288
rect 2652 25248 2688 25276
rect 2682 25236 2688 25248
rect 2740 25239 2752 25285
rect 2961 25279 3019 25285
rect 2961 25276 2973 25279
rect 2792 25248 2973 25276
rect 2740 25236 2746 25239
rect 2792 25220 2820 25248
rect 2961 25245 2973 25248
rect 3007 25245 3019 25279
rect 2961 25239 3019 25245
rect 4246 25236 4252 25288
rect 4304 25236 4310 25288
rect 5074 25276 5080 25288
rect 5035 25248 5080 25276
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 6914 25236 6920 25288
rect 6972 25276 6978 25288
rect 7009 25279 7067 25285
rect 7009 25276 7021 25279
rect 6972 25248 7021 25276
rect 6972 25236 6978 25248
rect 7009 25245 7021 25248
rect 7055 25245 7067 25279
rect 7742 25276 7748 25288
rect 7703 25248 7748 25276
rect 7009 25239 7067 25245
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 8389 25279 8447 25285
rect 8389 25245 8401 25279
rect 8435 25276 8447 25279
rect 8478 25276 8484 25288
rect 8435 25248 8484 25276
rect 8435 25245 8447 25248
rect 8389 25239 8447 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 9585 25279 9643 25285
rect 9585 25245 9597 25279
rect 9631 25276 9643 25279
rect 9784 25276 9812 25304
rect 9631 25248 9812 25276
rect 9631 25245 9643 25248
rect 9585 25239 9643 25245
rect 10318 25236 10324 25288
rect 10376 25276 10382 25288
rect 10413 25279 10471 25285
rect 10413 25276 10425 25279
rect 10376 25248 10425 25276
rect 10376 25236 10382 25248
rect 10413 25245 10425 25248
rect 10459 25245 10471 25279
rect 10520 25276 10548 25316
rect 10669 25279 10727 25285
rect 10669 25276 10681 25279
rect 10520 25248 10681 25276
rect 10413 25239 10471 25245
rect 10669 25245 10681 25248
rect 10715 25245 10727 25279
rect 12250 25276 12256 25288
rect 12211 25248 12256 25276
rect 10669 25239 10727 25245
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12526 25276 12532 25288
rect 12487 25248 12532 25276
rect 12526 25236 12532 25248
rect 12584 25236 12590 25288
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 12713 25279 12771 25285
rect 12713 25276 12725 25279
rect 12676 25248 12725 25276
rect 12676 25236 12682 25248
rect 12713 25245 12725 25248
rect 12759 25245 12771 25279
rect 13354 25276 13360 25288
rect 13315 25248 13360 25276
rect 12713 25239 12771 25245
rect 13354 25236 13360 25248
rect 13412 25236 13418 25288
rect 19426 25276 19432 25288
rect 19387 25248 19432 25276
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 20530 25236 20536 25288
rect 20588 25276 20594 25288
rect 22014 25279 22072 25285
rect 22014 25276 22026 25279
rect 20588 25248 22026 25276
rect 20588 25236 20594 25248
rect 22014 25245 22026 25248
rect 22060 25245 22072 25279
rect 22014 25239 22072 25245
rect 22281 25279 22339 25285
rect 22281 25245 22293 25279
rect 22327 25276 22339 25279
rect 22370 25276 22376 25288
rect 22327 25248 22376 25276
rect 22327 25245 22339 25248
rect 22281 25239 22339 25245
rect 22370 25236 22376 25248
rect 22428 25236 22434 25288
rect 2774 25168 2780 25220
rect 2832 25168 2838 25220
rect 3973 25211 4031 25217
rect 3973 25177 3985 25211
rect 4019 25208 4031 25211
rect 4062 25208 4068 25220
rect 4019 25180 4068 25208
rect 4019 25177 4031 25180
rect 3973 25171 4031 25177
rect 4062 25168 4068 25180
rect 4120 25168 4126 25220
rect 5626 25208 5632 25220
rect 4356 25180 5632 25208
rect 2130 25100 2136 25152
rect 2188 25140 2194 25152
rect 4356 25140 4384 25180
rect 5626 25168 5632 25180
rect 5684 25168 5690 25220
rect 9769 25211 9827 25217
rect 9769 25177 9781 25211
rect 9815 25208 9827 25211
rect 11054 25208 11060 25220
rect 9815 25180 11060 25208
rect 9815 25177 9827 25180
rect 9769 25171 9827 25177
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 12345 25211 12403 25217
rect 12345 25177 12357 25211
rect 12391 25208 12403 25211
rect 13446 25208 13452 25220
rect 12391 25180 13452 25208
rect 12391 25177 12403 25180
rect 12345 25171 12403 25177
rect 13446 25168 13452 25180
rect 13504 25168 13510 25220
rect 20441 25211 20499 25217
rect 20441 25177 20453 25211
rect 20487 25208 20499 25211
rect 21634 25208 21640 25220
rect 20487 25180 21640 25208
rect 20487 25177 20499 25180
rect 20441 25171 20499 25177
rect 20640 25152 20668 25180
rect 21634 25168 21640 25180
rect 21692 25168 21698 25220
rect 2188 25112 4384 25140
rect 4433 25143 4491 25149
rect 2188 25100 2194 25112
rect 4433 25109 4445 25143
rect 4479 25140 4491 25143
rect 4614 25140 4620 25152
rect 4479 25112 4620 25140
rect 4479 25109 4491 25112
rect 4433 25103 4491 25109
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 4890 25140 4896 25152
rect 4851 25112 4896 25140
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 9953 25143 10011 25149
rect 9953 25109 9965 25143
rect 9999 25140 10011 25143
rect 10594 25140 10600 25152
rect 9999 25112 10600 25140
rect 9999 25109 10011 25112
rect 9953 25103 10011 25109
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 10686 25100 10692 25152
rect 10744 25140 10750 25152
rect 11514 25140 11520 25152
rect 10744 25112 11520 25140
rect 10744 25100 10750 25112
rect 11514 25100 11520 25112
rect 11572 25140 11578 25152
rect 11793 25143 11851 25149
rect 11793 25140 11805 25143
rect 11572 25112 11805 25140
rect 11572 25100 11578 25112
rect 11793 25109 11805 25112
rect 11839 25109 11851 25143
rect 17770 25140 17776 25152
rect 17731 25112 17776 25140
rect 11793 25103 11851 25109
rect 17770 25100 17776 25112
rect 17828 25140 17834 25152
rect 18233 25143 18291 25149
rect 18233 25140 18245 25143
rect 17828 25112 18245 25140
rect 17828 25100 17834 25112
rect 18233 25109 18245 25112
rect 18279 25140 18291 25143
rect 18785 25143 18843 25149
rect 18785 25140 18797 25143
rect 18279 25112 18797 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 18785 25109 18797 25112
rect 18831 25109 18843 25143
rect 18785 25103 18843 25109
rect 19613 25143 19671 25149
rect 19613 25109 19625 25143
rect 19659 25140 19671 25143
rect 20070 25140 20076 25152
rect 19659 25112 20076 25140
rect 19659 25109 19671 25112
rect 19613 25103 19671 25109
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 20241 25143 20299 25149
rect 20241 25109 20253 25143
rect 20287 25140 20299 25143
rect 20530 25140 20536 25152
rect 20287 25112 20536 25140
rect 20287 25109 20299 25112
rect 20241 25103 20299 25109
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 20622 25100 20628 25152
rect 20680 25100 20686 25152
rect 1104 25050 22976 25072
rect 1104 24998 6378 25050
rect 6430 24998 6442 25050
rect 6494 24998 6506 25050
rect 6558 24998 6570 25050
rect 6622 24998 6634 25050
rect 6686 24998 11806 25050
rect 11858 24998 11870 25050
rect 11922 24998 11934 25050
rect 11986 24998 11998 25050
rect 12050 24998 12062 25050
rect 12114 24998 17234 25050
rect 17286 24998 17298 25050
rect 17350 24998 17362 25050
rect 17414 24998 17426 25050
rect 17478 24998 17490 25050
rect 17542 24998 22662 25050
rect 22714 24998 22726 25050
rect 22778 24998 22790 25050
rect 22842 24998 22854 25050
rect 22906 24998 22918 25050
rect 22970 24998 22976 25050
rect 1104 24976 22976 24998
rect 2038 24896 2044 24948
rect 2096 24936 2102 24948
rect 6178 24936 6184 24948
rect 2096 24908 6184 24936
rect 2096 24896 2102 24908
rect 6178 24896 6184 24908
rect 6236 24896 6242 24948
rect 8846 24896 8852 24948
rect 8904 24936 8910 24948
rect 9927 24939 9985 24945
rect 9927 24936 9939 24939
rect 8904 24908 9939 24936
rect 8904 24896 8910 24908
rect 9927 24905 9939 24908
rect 9973 24936 9985 24939
rect 9973 24908 10640 24936
rect 9973 24905 9985 24908
rect 9927 24899 9985 24905
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 2774 24868 2780 24880
rect 2372 24840 2780 24868
rect 2372 24828 2378 24840
rect 2774 24828 2780 24840
rect 2832 24868 2838 24880
rect 2832 24840 3004 24868
rect 2832 24828 2838 24840
rect 2682 24760 2688 24812
rect 2740 24809 2746 24812
rect 2976 24809 3004 24840
rect 3418 24828 3424 24880
rect 3476 24868 3482 24880
rect 3697 24871 3755 24877
rect 3697 24868 3709 24871
rect 3476 24840 3709 24868
rect 3476 24828 3482 24840
rect 3697 24837 3709 24840
rect 3743 24837 3755 24871
rect 3697 24831 3755 24837
rect 4798 24828 4804 24880
rect 4856 24868 4862 24880
rect 7098 24868 7104 24880
rect 4856 24840 7104 24868
rect 4856 24828 4862 24840
rect 7098 24828 7104 24840
rect 7156 24828 7162 24880
rect 10137 24871 10195 24877
rect 10137 24837 10149 24871
rect 10183 24868 10195 24871
rect 10502 24868 10508 24880
rect 10183 24840 10508 24868
rect 10183 24837 10195 24840
rect 10137 24831 10195 24837
rect 10502 24828 10508 24840
rect 10560 24828 10566 24880
rect 3602 24809 3608 24812
rect 2740 24800 2752 24809
rect 2961 24803 3019 24809
rect 2740 24772 2785 24800
rect 2740 24763 2752 24772
rect 2961 24769 2973 24803
rect 3007 24769 3019 24803
rect 2961 24763 3019 24769
rect 3581 24803 3608 24809
rect 3581 24769 3593 24803
rect 3581 24763 3608 24769
rect 2740 24760 2746 24763
rect 3602 24760 3608 24763
rect 3660 24760 3666 24812
rect 3789 24803 3847 24809
rect 3789 24798 3801 24803
rect 3712 24770 3801 24798
rect 3326 24692 3332 24744
rect 3384 24732 3390 24744
rect 3712 24732 3740 24770
rect 3789 24769 3801 24770
rect 3835 24769 3847 24803
rect 3789 24763 3847 24769
rect 3973 24803 4031 24809
rect 3973 24769 3985 24803
rect 4019 24769 4031 24803
rect 3973 24763 4031 24769
rect 3384 24704 3740 24732
rect 3384 24692 3390 24704
rect 3988 24664 4016 24763
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4893 24803 4951 24809
rect 4893 24800 4905 24803
rect 4120 24772 4905 24800
rect 4120 24760 4126 24772
rect 4893 24769 4905 24772
rect 4939 24800 4951 24803
rect 5074 24800 5080 24812
rect 4939 24772 5080 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5537 24803 5595 24809
rect 5537 24790 5549 24803
rect 5460 24769 5549 24790
rect 5583 24769 5595 24803
rect 5460 24763 5595 24769
rect 5460 24762 5580 24763
rect 4982 24692 4988 24744
rect 5040 24732 5046 24744
rect 5460 24732 5488 24762
rect 6270 24760 6276 24812
rect 6328 24800 6334 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6328 24772 6561 24800
rect 6328 24760 6334 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24800 7435 24803
rect 7466 24800 7472 24812
rect 7423 24772 7472 24800
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 7558 24760 7564 24812
rect 7616 24800 7622 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 7616 24772 7849 24800
rect 7616 24760 7622 24772
rect 7837 24769 7849 24772
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8352 24772 8493 24800
rect 8352 24760 8358 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24769 9183 24803
rect 10612 24800 10640 24908
rect 10962 24896 10968 24948
rect 11020 24936 11026 24948
rect 12621 24939 12679 24945
rect 12621 24936 12633 24939
rect 11020 24908 12633 24936
rect 11020 24896 11026 24908
rect 12621 24905 12633 24908
rect 12667 24905 12679 24939
rect 12621 24899 12679 24905
rect 20073 24939 20131 24945
rect 20073 24905 20085 24939
rect 20119 24936 20131 24939
rect 21082 24936 21088 24948
rect 20119 24908 21088 24936
rect 20119 24905 20131 24908
rect 20073 24899 20131 24905
rect 10781 24871 10839 24877
rect 10781 24837 10793 24871
rect 10827 24868 10839 24871
rect 14274 24868 14280 24880
rect 10827 24840 11284 24868
rect 10827 24837 10839 24840
rect 10781 24831 10839 24837
rect 11149 24803 11207 24809
rect 11149 24800 11161 24803
rect 10612 24772 11161 24800
rect 9125 24763 9183 24769
rect 11149 24769 11161 24772
rect 11195 24769 11207 24803
rect 11149 24763 11207 24769
rect 5040 24704 5488 24732
rect 9140 24732 9168 24763
rect 9140 24704 10640 24732
rect 5040 24692 5046 24704
rect 5258 24664 5264 24676
rect 3988 24636 5264 24664
rect 4264 24608 4292 24636
rect 5258 24624 5264 24636
rect 5316 24624 5322 24676
rect 5350 24624 5356 24676
rect 5408 24664 5414 24676
rect 9309 24667 9367 24673
rect 5408 24636 5453 24664
rect 5408 24624 5414 24636
rect 9309 24633 9321 24667
rect 9355 24664 9367 24667
rect 9674 24664 9680 24676
rect 9355 24636 9680 24664
rect 9355 24633 9367 24636
rect 9309 24627 9367 24633
rect 9674 24624 9680 24636
rect 9732 24624 9738 24676
rect 9769 24667 9827 24673
rect 9769 24633 9781 24667
rect 9815 24664 9827 24667
rect 9858 24664 9864 24676
rect 9815 24636 9864 24664
rect 9815 24633 9827 24636
rect 9769 24627 9827 24633
rect 9858 24624 9864 24636
rect 9916 24624 9922 24676
rect 10612 24673 10640 24704
rect 10686 24692 10692 24744
rect 10744 24732 10750 24744
rect 11256 24732 11284 24840
rect 12406 24840 14280 24868
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11664 24772 11713 24800
rect 11664 24760 11670 24772
rect 11701 24769 11713 24772
rect 11747 24800 11759 24803
rect 12406 24800 12434 24840
rect 14274 24828 14280 24840
rect 14332 24828 14338 24880
rect 19334 24828 19340 24880
rect 19392 24828 19398 24880
rect 19437 24871 19495 24877
rect 19437 24837 19449 24871
rect 19483 24868 19495 24871
rect 19483 24840 19564 24868
rect 19483 24837 19495 24840
rect 19437 24831 19495 24837
rect 12802 24800 12808 24812
rect 11747 24772 12434 24800
rect 12763 24772 12808 24800
rect 11747 24769 11759 24772
rect 11701 24763 11759 24769
rect 12802 24760 12808 24772
rect 12860 24760 12866 24812
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 18601 24803 18659 24809
rect 18601 24800 18613 24803
rect 17460 24772 18613 24800
rect 17460 24760 17466 24772
rect 18601 24769 18613 24772
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19352 24800 19380 24828
rect 19291 24772 19380 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 12161 24735 12219 24741
rect 10744 24704 12020 24732
rect 10744 24692 10750 24704
rect 11992 24673 12020 24704
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 17034 24732 17040 24744
rect 12207 24704 17040 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 19536 24732 19564 24840
rect 20088 24732 20116 24899
rect 21082 24896 21088 24908
rect 21140 24936 21146 24948
rect 21634 24936 21640 24948
rect 21140 24908 21640 24936
rect 21140 24896 21146 24908
rect 21634 24896 21640 24908
rect 21692 24896 21698 24948
rect 20162 24828 20168 24880
rect 20220 24868 20226 24880
rect 20990 24868 20996 24880
rect 20220 24840 20996 24868
rect 20220 24828 20226 24840
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 21197 24803 21255 24809
rect 21197 24769 21209 24803
rect 21243 24800 21255 24803
rect 21542 24800 21548 24812
rect 21243 24772 21548 24800
rect 21243 24769 21255 24772
rect 21197 24763 21255 24769
rect 21542 24760 21548 24772
rect 21600 24760 21606 24812
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 22152 24772 22201 24800
rect 22152 24760 22158 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 18104 24704 20116 24732
rect 21453 24735 21511 24741
rect 18104 24692 18110 24704
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22370 24732 22376 24744
rect 21499 24704 22376 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 22370 24692 22376 24704
rect 22428 24692 22434 24744
rect 10597 24667 10655 24673
rect 10597 24633 10609 24667
rect 10643 24633 10655 24667
rect 10597 24627 10655 24633
rect 11977 24667 12035 24673
rect 11977 24633 11989 24667
rect 12023 24633 12035 24667
rect 11977 24627 12035 24633
rect 18141 24667 18199 24673
rect 18141 24633 18153 24667
rect 18187 24664 18199 24667
rect 19794 24664 19800 24676
rect 18187 24636 19800 24664
rect 18187 24633 18199 24636
rect 18141 24627 18199 24633
rect 19794 24624 19800 24636
rect 19852 24624 19858 24676
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2774 24556 2780 24608
rect 2832 24596 2838 24608
rect 3421 24599 3479 24605
rect 3421 24596 3433 24599
rect 2832 24568 3433 24596
rect 2832 24556 2838 24568
rect 3421 24565 3433 24568
rect 3467 24565 3479 24599
rect 3421 24559 3479 24565
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 4154 24596 4160 24608
rect 3660 24568 4160 24596
rect 3660 24556 3666 24568
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 4246 24556 4252 24608
rect 4304 24556 4310 24608
rect 4338 24556 4344 24608
rect 4396 24596 4402 24608
rect 4433 24599 4491 24605
rect 4433 24596 4445 24599
rect 4396 24568 4445 24596
rect 4396 24556 4402 24568
rect 4433 24565 4445 24568
rect 4479 24565 4491 24599
rect 4433 24559 4491 24565
rect 4522 24556 4528 24608
rect 4580 24596 4586 24608
rect 4617 24599 4675 24605
rect 4617 24596 4629 24599
rect 4580 24568 4629 24596
rect 4580 24556 4586 24568
rect 4617 24565 4629 24568
rect 4663 24565 4675 24599
rect 4617 24559 4675 24565
rect 5074 24556 5080 24608
rect 5132 24596 5138 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 5132 24568 7205 24596
rect 5132 24556 5138 24568
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 8570 24596 8576 24608
rect 8531 24568 8576 24596
rect 7193 24559 7251 24565
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 9950 24596 9956 24608
rect 9863 24568 9956 24596
rect 9950 24556 9956 24568
rect 10008 24596 10014 24608
rect 10502 24596 10508 24608
rect 10008 24568 10508 24596
rect 10008 24556 10014 24568
rect 10502 24556 10508 24568
rect 10560 24556 10566 24608
rect 10686 24556 10692 24608
rect 10744 24596 10750 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10744 24568 10793 24596
rect 10744 24556 10750 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 17497 24599 17555 24605
rect 17497 24565 17509 24599
rect 17543 24596 17555 24599
rect 17770 24596 17776 24608
rect 17543 24568 17776 24596
rect 17543 24565 17555 24568
rect 17497 24559 17555 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18690 24596 18696 24608
rect 18651 24568 18696 24596
rect 18690 24556 18696 24568
rect 18748 24556 18754 24608
rect 19610 24596 19616 24608
rect 19571 24568 19616 24596
rect 19610 24556 19616 24568
rect 19668 24556 19674 24608
rect 21450 24556 21456 24608
rect 21508 24596 21514 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21508 24568 22017 24596
rect 21508 24556 21514 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22005 24559 22063 24565
rect 1104 24506 22816 24528
rect 1104 24454 3664 24506
rect 3716 24454 3728 24506
rect 3780 24454 3792 24506
rect 3844 24454 3856 24506
rect 3908 24454 3920 24506
rect 3972 24454 9092 24506
rect 9144 24454 9156 24506
rect 9208 24454 9220 24506
rect 9272 24454 9284 24506
rect 9336 24454 9348 24506
rect 9400 24454 14520 24506
rect 14572 24454 14584 24506
rect 14636 24454 14648 24506
rect 14700 24454 14712 24506
rect 14764 24454 14776 24506
rect 14828 24454 19948 24506
rect 20000 24454 20012 24506
rect 20064 24454 20076 24506
rect 20128 24454 20140 24506
rect 20192 24454 20204 24506
rect 20256 24454 22816 24506
rect 1104 24432 22816 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 4246 24392 4252 24404
rect 1728 24364 4252 24392
rect 1728 24352 1734 24364
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 4430 24352 4436 24404
rect 4488 24392 4494 24404
rect 5169 24395 5227 24401
rect 5169 24392 5181 24395
rect 4488 24364 5181 24392
rect 4488 24352 4494 24364
rect 5169 24361 5181 24364
rect 5215 24361 5227 24395
rect 5169 24355 5227 24361
rect 4985 24327 5043 24333
rect 4985 24293 4997 24327
rect 5031 24293 5043 24327
rect 5184 24324 5212 24355
rect 5442 24352 5448 24404
rect 5500 24392 5506 24404
rect 8481 24395 8539 24401
rect 8481 24392 8493 24395
rect 5500 24364 8493 24392
rect 5500 24352 5506 24364
rect 8481 24361 8493 24364
rect 8527 24361 8539 24395
rect 9582 24392 9588 24404
rect 9543 24364 9588 24392
rect 8481 24355 8539 24361
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 10410 24392 10416 24404
rect 10371 24364 10416 24392
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 11146 24352 11152 24404
rect 11204 24392 11210 24404
rect 11701 24395 11759 24401
rect 11701 24392 11713 24395
rect 11204 24364 11713 24392
rect 11204 24352 11210 24364
rect 11701 24361 11713 24364
rect 11747 24361 11759 24395
rect 17402 24392 17408 24404
rect 17363 24364 17408 24392
rect 11701 24355 11759 24361
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 17586 24352 17592 24404
rect 17644 24392 17650 24404
rect 18693 24395 18751 24401
rect 18693 24392 18705 24395
rect 17644 24364 18705 24392
rect 17644 24352 17650 24364
rect 18693 24361 18705 24364
rect 18739 24361 18751 24395
rect 18693 24355 18751 24361
rect 18877 24395 18935 24401
rect 18877 24361 18889 24395
rect 18923 24392 18935 24395
rect 19426 24392 19432 24404
rect 18923 24364 19432 24392
rect 18923 24361 18935 24364
rect 18877 24355 18935 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 20073 24395 20131 24401
rect 20073 24392 20085 24395
rect 19668 24364 20085 24392
rect 19668 24352 19674 24364
rect 20073 24361 20085 24364
rect 20119 24361 20131 24395
rect 20073 24355 20131 24361
rect 20714 24352 20720 24404
rect 20772 24392 20778 24404
rect 20901 24395 20959 24401
rect 20901 24392 20913 24395
rect 20772 24364 20913 24392
rect 20772 24352 20778 24364
rect 20901 24361 20913 24364
rect 20947 24392 20959 24395
rect 21910 24392 21916 24404
rect 20947 24364 21916 24392
rect 20947 24361 20959 24364
rect 20901 24355 20959 24361
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 6638 24324 6644 24336
rect 5184 24296 5580 24324
rect 6599 24296 6644 24324
rect 4985 24287 5043 24293
rect 4433 24259 4491 24265
rect 4433 24225 4445 24259
rect 4479 24256 4491 24259
rect 4706 24256 4712 24268
rect 4479 24228 4712 24256
rect 4479 24225 4491 24228
rect 4433 24219 4491 24225
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 5000 24256 5028 24287
rect 5442 24256 5448 24268
rect 5000 24228 5448 24256
rect 5442 24216 5448 24228
rect 5500 24216 5506 24268
rect 2682 24148 2688 24200
rect 2740 24197 2746 24200
rect 2740 24188 2752 24197
rect 2961 24191 3019 24197
rect 2740 24160 2785 24188
rect 2740 24151 2752 24160
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3602 24188 3608 24200
rect 3007 24160 3608 24188
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 2740 24148 2746 24151
rect 2314 24080 2320 24132
rect 2372 24120 2378 24132
rect 2976 24120 3004 24151
rect 3602 24148 3608 24160
rect 3660 24148 3666 24200
rect 4154 24188 4160 24200
rect 4115 24160 4160 24188
rect 4154 24148 4160 24160
rect 4212 24148 4218 24200
rect 4249 24191 4307 24197
rect 4249 24157 4261 24191
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24188 4583 24191
rect 5074 24188 5080 24200
rect 4571 24184 4660 24188
rect 4816 24184 5080 24188
rect 4571 24160 5080 24184
rect 4571 24157 4583 24160
rect 4525 24151 4583 24157
rect 4632 24156 4844 24160
rect 2372 24092 3004 24120
rect 2372 24080 2378 24092
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 4264 24120 4292 24151
rect 5074 24148 5080 24160
rect 5132 24148 5138 24200
rect 4430 24120 4436 24132
rect 3476 24092 4436 24120
rect 3476 24080 3482 24092
rect 4430 24080 4436 24092
rect 4488 24080 4494 24132
rect 5350 24120 5356 24132
rect 5311 24092 5356 24120
rect 5350 24080 5356 24092
rect 5408 24080 5414 24132
rect 5552 24120 5580 24296
rect 6638 24284 6644 24296
rect 6696 24284 6702 24336
rect 7190 24284 7196 24336
rect 7248 24324 7254 24336
rect 7285 24327 7343 24333
rect 7285 24324 7297 24327
rect 7248 24296 7297 24324
rect 7248 24284 7254 24296
rect 7285 24293 7297 24296
rect 7331 24293 7343 24327
rect 7285 24287 7343 24293
rect 7466 24284 7472 24336
rect 7524 24324 7530 24336
rect 7929 24327 7987 24333
rect 7929 24324 7941 24327
rect 7524 24296 7941 24324
rect 7524 24284 7530 24296
rect 7929 24293 7941 24296
rect 7975 24293 7987 24327
rect 7929 24287 7987 24293
rect 8570 24284 8576 24336
rect 8628 24324 8634 24336
rect 13170 24324 13176 24336
rect 8628 24296 13176 24324
rect 8628 24284 8634 24296
rect 13170 24284 13176 24296
rect 13228 24284 13234 24336
rect 20441 24327 20499 24333
rect 20441 24293 20453 24327
rect 20487 24324 20499 24327
rect 21266 24324 21272 24336
rect 20487 24296 21272 24324
rect 20487 24293 20499 24296
rect 20441 24287 20499 24293
rect 21266 24284 21272 24296
rect 21324 24284 21330 24336
rect 10042 24216 10048 24268
rect 10100 24256 10106 24268
rect 10873 24259 10931 24265
rect 10873 24256 10885 24259
rect 10100 24228 10885 24256
rect 10100 24216 10106 24228
rect 10873 24225 10885 24228
rect 10919 24225 10931 24259
rect 10873 24219 10931 24225
rect 12342 24216 12348 24268
rect 12400 24256 12406 24268
rect 12437 24259 12495 24265
rect 12437 24256 12449 24259
rect 12400 24228 12449 24256
rect 12400 24216 12406 24228
rect 12437 24225 12449 24228
rect 12483 24225 12495 24259
rect 19334 24256 19340 24268
rect 12437 24219 12495 24225
rect 17236 24228 19340 24256
rect 5626 24148 5632 24200
rect 5684 24188 5690 24200
rect 6825 24191 6883 24197
rect 6825 24188 6837 24191
rect 5684 24160 6837 24188
rect 5684 24148 5690 24160
rect 6825 24157 6837 24160
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 9490 24148 9496 24200
rect 9548 24188 9554 24200
rect 10229 24191 10287 24197
rect 10229 24188 10241 24191
rect 9548 24160 10241 24188
rect 9548 24148 9554 24160
rect 10229 24157 10241 24160
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 11330 24188 11336 24200
rect 11287 24160 11336 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 17236 24197 17264 24228
rect 19334 24216 19340 24228
rect 19392 24216 19398 24268
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24188 16819 24191
rect 17221 24191 17279 24197
rect 17221 24188 17233 24191
rect 16807 24160 17233 24188
rect 16807 24157 16819 24160
rect 16761 24151 16819 24157
rect 17221 24157 17233 24160
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17678 24148 17684 24200
rect 17736 24188 17742 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 17736 24160 17877 24188
rect 17736 24148 17742 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 19058 24188 19064 24200
rect 18095 24160 19064 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 5998 24123 6056 24129
rect 5998 24120 6010 24123
rect 5552 24092 6010 24120
rect 5998 24089 6010 24092
rect 6044 24089 6056 24123
rect 6178 24120 6184 24132
rect 6139 24092 6184 24120
rect 5998 24083 6056 24089
rect 6178 24080 6184 24092
rect 6236 24080 6242 24132
rect 11057 24123 11115 24129
rect 11057 24089 11069 24123
rect 11103 24120 11115 24123
rect 11422 24120 11428 24132
rect 11103 24092 11428 24120
rect 11103 24089 11115 24092
rect 11057 24083 11115 24089
rect 11422 24080 11428 24092
rect 11480 24080 11486 24132
rect 18064 24120 18092 24151
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19242 24148 19248 24200
rect 19300 24188 19306 24200
rect 19610 24188 19616 24200
rect 19300 24160 19616 24188
rect 19300 24148 19306 24160
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 19978 24188 19984 24200
rect 19812 24160 19984 24188
rect 17880 24092 18092 24120
rect 18509 24123 18567 24129
rect 17880 24064 17908 24092
rect 18509 24089 18521 24123
rect 18555 24120 18567 24123
rect 19812 24120 19840 24160
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 22002 24188 22008 24200
rect 22060 24197 22066 24200
rect 21972 24160 22008 24188
rect 22002 24148 22008 24160
rect 22060 24151 22072 24197
rect 22281 24191 22339 24197
rect 22281 24157 22293 24191
rect 22327 24188 22339 24191
rect 22370 24188 22376 24200
rect 22327 24160 22376 24188
rect 22327 24157 22339 24160
rect 22281 24151 22339 24157
rect 22060 24148 22066 24151
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 22186 24120 22192 24132
rect 18555 24092 19840 24120
rect 19904 24092 21956 24120
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 1670 24052 1676 24064
rect 1627 24024 1676 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 5166 24061 5172 24064
rect 3973 24055 4031 24061
rect 3973 24052 3985 24055
rect 2556 24024 3985 24052
rect 2556 24012 2562 24024
rect 3973 24021 3985 24024
rect 4019 24021 4031 24055
rect 3973 24015 4031 24021
rect 5153 24055 5172 24061
rect 5153 24021 5165 24055
rect 5153 24015 5172 24021
rect 5166 24012 5172 24015
rect 5224 24012 5230 24064
rect 5810 24052 5816 24064
rect 5771 24024 5816 24052
rect 5810 24012 5816 24024
rect 5868 24012 5874 24064
rect 17862 24012 17868 24064
rect 17920 24012 17926 24064
rect 19904 24061 19932 24092
rect 18049 24055 18107 24061
rect 18049 24021 18061 24055
rect 18095 24052 18107 24055
rect 18709 24055 18767 24061
rect 18709 24052 18721 24055
rect 18095 24024 18721 24052
rect 18095 24021 18107 24024
rect 18049 24015 18107 24021
rect 18709 24021 18721 24024
rect 18755 24021 18767 24055
rect 18709 24015 18767 24021
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24021 19947 24055
rect 19889 24015 19947 24021
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 20073 24055 20131 24061
rect 20073 24052 20085 24055
rect 20036 24024 20085 24052
rect 20036 24012 20042 24024
rect 20073 24021 20085 24024
rect 20119 24021 20131 24055
rect 21928 24052 21956 24092
rect 22066 24092 22192 24120
rect 22066 24052 22094 24092
rect 22186 24080 22192 24092
rect 22244 24080 22250 24132
rect 21928 24024 22094 24052
rect 20073 24015 20131 24021
rect 1104 23962 22976 23984
rect 1104 23910 6378 23962
rect 6430 23910 6442 23962
rect 6494 23910 6506 23962
rect 6558 23910 6570 23962
rect 6622 23910 6634 23962
rect 6686 23910 11806 23962
rect 11858 23910 11870 23962
rect 11922 23910 11934 23962
rect 11986 23910 11998 23962
rect 12050 23910 12062 23962
rect 12114 23910 17234 23962
rect 17286 23910 17298 23962
rect 17350 23910 17362 23962
rect 17414 23910 17426 23962
rect 17478 23910 17490 23962
rect 17542 23910 22662 23962
rect 22714 23910 22726 23962
rect 22778 23910 22790 23962
rect 22842 23910 22854 23962
rect 22906 23910 22918 23962
rect 22970 23910 22976 23962
rect 1104 23888 22976 23910
rect 3142 23808 3148 23860
rect 3200 23848 3206 23860
rect 3881 23851 3939 23857
rect 3881 23848 3893 23851
rect 3200 23820 3893 23848
rect 3200 23808 3206 23820
rect 3881 23817 3893 23820
rect 3927 23848 3939 23851
rect 4062 23848 4068 23860
rect 3927 23820 4068 23848
rect 3927 23817 3939 23820
rect 3881 23811 3939 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 4212 23820 5825 23848
rect 4212 23808 4218 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 6178 23808 6184 23860
rect 6236 23848 6242 23860
rect 6549 23851 6607 23857
rect 6549 23848 6561 23851
rect 6236 23820 6561 23848
rect 6236 23808 6242 23820
rect 6549 23817 6561 23820
rect 6595 23817 6607 23851
rect 6549 23811 6607 23817
rect 10870 23808 10876 23860
rect 10928 23848 10934 23860
rect 10965 23851 11023 23857
rect 10965 23848 10977 23851
rect 10928 23820 10977 23848
rect 10928 23808 10934 23820
rect 10965 23817 10977 23820
rect 11011 23817 11023 23851
rect 17586 23848 17592 23860
rect 17547 23820 17592 23848
rect 10965 23811 11023 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 19334 23848 19340 23860
rect 18340 23820 19340 23848
rect 4706 23780 4712 23792
rect 3436 23752 4712 23780
rect 1578 23712 1584 23724
rect 1539 23684 1584 23712
rect 1578 23672 1584 23684
rect 1636 23672 1642 23724
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23712 2191 23715
rect 2222 23712 2228 23724
rect 2179 23684 2228 23712
rect 2179 23681 2191 23684
rect 2133 23675 2191 23681
rect 2222 23672 2228 23684
rect 2280 23672 2286 23724
rect 2498 23712 2504 23724
rect 2459 23684 2504 23712
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 3436 23721 3464 23752
rect 4706 23740 4712 23752
rect 4764 23740 4770 23792
rect 5074 23740 5080 23792
rect 5132 23740 5138 23792
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 8110 23780 8116 23792
rect 5408 23752 6868 23780
rect 8023 23752 8116 23780
rect 5408 23740 5414 23752
rect 3053 23715 3111 23721
rect 3053 23681 3065 23715
rect 3099 23712 3111 23715
rect 3421 23715 3479 23721
rect 3099 23684 3372 23712
rect 3099 23681 3111 23684
rect 3053 23675 3111 23681
rect 2590 23644 2596 23656
rect 2551 23616 2596 23644
rect 2590 23604 2596 23616
rect 2648 23604 2654 23656
rect 3142 23468 3148 23520
rect 3200 23508 3206 23520
rect 3344 23508 3372 23684
rect 3421 23681 3433 23715
rect 3467 23681 3479 23715
rect 3421 23675 3479 23681
rect 4430 23672 4436 23724
rect 4488 23712 4494 23724
rect 4994 23715 5052 23721
rect 4994 23712 5006 23715
rect 4488 23684 5006 23712
rect 4488 23672 4494 23684
rect 4994 23681 5006 23684
rect 5040 23681 5052 23715
rect 5092 23712 5120 23740
rect 5092 23684 5396 23712
rect 4994 23675 5052 23681
rect 5368 23656 5396 23684
rect 5902 23672 5908 23724
rect 5960 23712 5966 23724
rect 6730 23712 6736 23724
rect 5960 23684 6005 23712
rect 6691 23684 6736 23712
rect 5960 23672 5966 23684
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 6840 23721 6868 23752
rect 8110 23740 8116 23752
rect 8168 23780 8174 23792
rect 12342 23780 12348 23792
rect 8168 23752 12348 23780
rect 8168 23740 8174 23752
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 16666 23740 16672 23792
rect 16724 23780 16730 23792
rect 17405 23783 17463 23789
rect 17405 23780 17417 23783
rect 16724 23752 17417 23780
rect 16724 23740 16730 23752
rect 17405 23749 17417 23752
rect 17451 23780 17463 23783
rect 17862 23780 17868 23792
rect 17451 23752 17868 23780
rect 17451 23749 17463 23752
rect 17405 23743 17463 23749
rect 17862 23740 17868 23752
rect 17920 23740 17926 23792
rect 18340 23789 18368 23820
rect 19334 23808 19340 23820
rect 19392 23848 19398 23860
rect 20438 23848 20444 23860
rect 19392 23820 20444 23848
rect 19392 23808 19398 23820
rect 20438 23808 20444 23820
rect 20496 23848 20502 23860
rect 20714 23848 20720 23860
rect 20496 23820 20720 23848
rect 20496 23808 20502 23820
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 22005 23851 22063 23857
rect 22005 23817 22017 23851
rect 22051 23817 22063 23851
rect 22005 23811 22063 23817
rect 18325 23783 18383 23789
rect 18325 23749 18337 23783
rect 18371 23749 18383 23783
rect 21208 23783 21266 23789
rect 18325 23743 18383 23749
rect 18432 23752 19472 23780
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7561 23675 7619 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23712 11207 23715
rect 11238 23712 11244 23724
rect 11195 23684 11244 23712
rect 11195 23681 11207 23684
rect 11149 23675 11207 23681
rect 5258 23644 5264 23656
rect 5219 23616 5264 23644
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 5350 23604 5356 23656
rect 5408 23644 5414 23656
rect 7392 23644 7420 23675
rect 5408 23616 7420 23644
rect 5408 23604 5414 23616
rect 5442 23536 5448 23588
rect 5500 23576 5506 23588
rect 7576 23576 7604 23675
rect 11238 23672 11244 23684
rect 11296 23672 11302 23724
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 18046 23712 18052 23724
rect 18007 23684 18052 23712
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 18432 23721 18460 23752
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23681 18475 23715
rect 19058 23712 19064 23724
rect 19019 23684 19064 23712
rect 18417 23675 18475 23681
rect 5500 23548 7604 23576
rect 18248 23576 18276 23675
rect 19058 23672 19064 23684
rect 19116 23672 19122 23724
rect 19334 23712 19340 23724
rect 19295 23684 19340 23712
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 19444 23721 19472 23752
rect 21208 23749 21220 23783
rect 21254 23780 21266 23783
rect 22020 23780 22048 23811
rect 21254 23752 22048 23780
rect 21254 23749 21266 23752
rect 21208 23743 21266 23749
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23712 19487 23715
rect 19518 23712 19524 23724
rect 19475 23684 19524 23712
rect 19475 23681 19487 23684
rect 19429 23675 19487 23681
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 21358 23712 21364 23724
rect 20456 23684 21364 23712
rect 19153 23647 19211 23653
rect 19153 23613 19165 23647
rect 19199 23644 19211 23647
rect 20456 23644 20484 23684
rect 21358 23672 21364 23684
rect 21416 23672 21422 23724
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 19199 23616 20484 23644
rect 21453 23647 21511 23653
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 21453 23613 21465 23647
rect 21499 23644 21511 23647
rect 21542 23644 21548 23656
rect 21499 23616 21548 23644
rect 21499 23613 21511 23616
rect 21453 23607 21511 23613
rect 21542 23604 21548 23616
rect 21600 23644 21606 23656
rect 22370 23644 22376 23656
rect 21600 23616 22376 23644
rect 21600 23604 21606 23616
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 19426 23576 19432 23588
rect 18248 23548 19432 23576
rect 5500 23536 5506 23548
rect 19426 23536 19432 23548
rect 19484 23536 19490 23588
rect 19613 23579 19671 23585
rect 19613 23545 19625 23579
rect 19659 23576 19671 23579
rect 19659 23548 20576 23576
rect 19659 23545 19671 23548
rect 19613 23539 19671 23545
rect 5350 23508 5356 23520
rect 3200 23480 5356 23508
rect 3200 23468 3206 23480
rect 5350 23468 5356 23480
rect 5408 23468 5414 23520
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 7469 23511 7527 23517
rect 7469 23508 7481 23511
rect 6880 23480 7481 23508
rect 6880 23468 6886 23480
rect 7469 23477 7481 23480
rect 7515 23477 7527 23511
rect 18598 23508 18604 23520
rect 18559 23480 18604 23508
rect 7469 23471 7527 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 20073 23511 20131 23517
rect 20073 23477 20085 23511
rect 20119 23508 20131 23511
rect 20438 23508 20444 23520
rect 20119 23480 20444 23508
rect 20119 23477 20131 23480
rect 20073 23471 20131 23477
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 20548 23508 20576 23548
rect 21266 23508 21272 23520
rect 20548 23480 21272 23508
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 1104 23418 22816 23440
rect 1104 23366 3664 23418
rect 3716 23366 3728 23418
rect 3780 23366 3792 23418
rect 3844 23366 3856 23418
rect 3908 23366 3920 23418
rect 3972 23366 9092 23418
rect 9144 23366 9156 23418
rect 9208 23366 9220 23418
rect 9272 23366 9284 23418
rect 9336 23366 9348 23418
rect 9400 23366 14520 23418
rect 14572 23366 14584 23418
rect 14636 23366 14648 23418
rect 14700 23366 14712 23418
rect 14764 23366 14776 23418
rect 14828 23366 19948 23418
rect 20000 23366 20012 23418
rect 20064 23366 20076 23418
rect 20128 23366 20140 23418
rect 20192 23366 20204 23418
rect 20256 23366 22816 23418
rect 1104 23344 22816 23366
rect 2961 23307 3019 23313
rect 2961 23273 2973 23307
rect 3007 23304 3019 23307
rect 3418 23304 3424 23316
rect 3007 23276 3424 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 5902 23304 5908 23316
rect 5863 23276 5908 23304
rect 5902 23264 5908 23276
rect 5960 23264 5966 23316
rect 6086 23264 6092 23316
rect 6144 23304 6150 23316
rect 7745 23307 7803 23313
rect 7745 23304 7757 23307
rect 6144 23276 7757 23304
rect 6144 23264 6150 23276
rect 7745 23273 7757 23276
rect 7791 23304 7803 23307
rect 9858 23304 9864 23316
rect 7791 23276 9864 23304
rect 7791 23273 7803 23276
rect 7745 23267 7803 23273
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 16850 23304 16856 23316
rect 16811 23276 16856 23304
rect 16850 23264 16856 23276
rect 16908 23304 16914 23316
rect 16908 23276 18736 23304
rect 16908 23264 16914 23276
rect 4890 23236 4896 23248
rect 2746 23208 4896 23236
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 1848 23103 1906 23109
rect 1848 23069 1860 23103
rect 1894 23100 1906 23103
rect 2746 23100 2774 23208
rect 4890 23196 4896 23208
rect 4948 23196 4954 23248
rect 6914 23196 6920 23248
rect 6972 23236 6978 23248
rect 7193 23239 7251 23245
rect 7193 23236 7205 23239
rect 6972 23208 7205 23236
rect 6972 23196 6978 23208
rect 7193 23205 7205 23208
rect 7239 23205 7251 23239
rect 17034 23236 17040 23248
rect 16995 23208 17040 23236
rect 7193 23199 7251 23205
rect 17034 23196 17040 23208
rect 17092 23196 17098 23248
rect 17862 23236 17868 23248
rect 17823 23208 17868 23236
rect 17862 23196 17868 23208
rect 17920 23196 17926 23248
rect 18708 23245 18736 23276
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 19484 23276 19809 23304
rect 19484 23264 19490 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 19797 23267 19855 23273
rect 19981 23307 20039 23313
rect 19981 23273 19993 23307
rect 20027 23304 20039 23307
rect 20346 23304 20352 23316
rect 20027 23276 20352 23304
rect 20027 23273 20039 23276
rect 19981 23267 20039 23273
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 20898 23264 20904 23316
rect 20956 23304 20962 23316
rect 20956 23276 22232 23304
rect 20956 23264 20962 23276
rect 18693 23239 18751 23245
rect 18693 23205 18705 23239
rect 18739 23205 18751 23239
rect 18693 23199 18751 23205
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 22094 23236 22100 23248
rect 18923 23208 22100 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 22094 23196 22100 23208
rect 22152 23196 22158 23248
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 5350 23168 5356 23180
rect 3016 23140 4476 23168
rect 3016 23128 3022 23140
rect 1894 23072 2774 23100
rect 1894 23069 1906 23072
rect 1848 23063 1906 23069
rect 2866 23060 2872 23112
rect 2924 23100 2930 23112
rect 3142 23100 3148 23112
rect 2924 23072 3148 23100
rect 2924 23060 2930 23072
rect 3142 23060 3148 23072
rect 3200 23060 3206 23112
rect 4154 23109 4160 23112
rect 4152 23100 4160 23109
rect 4115 23072 4160 23100
rect 4152 23063 4160 23072
rect 4154 23060 4160 23063
rect 4212 23060 4218 23112
rect 4448 23109 4476 23140
rect 5276 23140 5356 23168
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4448 23103 4527 23109
rect 4448 23072 4481 23103
rect 4341 23063 4399 23069
rect 4469 23069 4481 23072
rect 4515 23069 4527 23103
rect 4469 23063 4527 23069
rect 2958 22992 2964 23044
rect 3016 23032 3022 23044
rect 4062 23032 4068 23044
rect 3016 23004 4068 23032
rect 3016 22992 3022 23004
rect 4062 22992 4068 23004
rect 4120 23032 4126 23044
rect 4249 23035 4307 23041
rect 4249 23032 4261 23035
rect 4120 23004 4261 23032
rect 4120 22992 4126 23004
rect 4249 23001 4261 23004
rect 4295 23001 4307 23035
rect 4356 23032 4384 23063
rect 4614 23060 4620 23112
rect 4672 23100 4678 23112
rect 5276 23109 5304 23140
rect 5350 23128 5356 23140
rect 5408 23128 5414 23180
rect 18230 23128 18236 23180
rect 18288 23168 18294 23180
rect 18417 23171 18475 23177
rect 18417 23168 18429 23171
rect 18288 23140 18429 23168
rect 18288 23128 18294 23140
rect 18417 23137 18429 23140
rect 18463 23168 18475 23171
rect 20070 23168 20076 23180
rect 18463 23140 20076 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 20070 23128 20076 23140
rect 20128 23168 20134 23180
rect 20622 23168 20628 23180
rect 20128 23140 20628 23168
rect 20128 23128 20134 23140
rect 20622 23128 20628 23140
rect 20680 23128 20686 23180
rect 21082 23128 21088 23180
rect 21140 23168 21146 23180
rect 21177 23171 21235 23177
rect 21177 23168 21189 23171
rect 21140 23140 21189 23168
rect 21140 23128 21146 23140
rect 21177 23137 21189 23140
rect 21223 23137 21235 23171
rect 21177 23131 21235 23137
rect 21358 23128 21364 23180
rect 21416 23168 21422 23180
rect 21637 23171 21695 23177
rect 21637 23168 21649 23171
rect 21416 23140 21649 23168
rect 21416 23128 21422 23140
rect 21637 23137 21649 23140
rect 21683 23137 21695 23171
rect 21637 23131 21695 23137
rect 5261 23103 5319 23109
rect 4672 23072 4717 23100
rect 4672 23060 4678 23072
rect 5261 23069 5273 23103
rect 5307 23069 5319 23103
rect 6086 23100 6092 23112
rect 6047 23072 6092 23100
rect 5261 23063 5319 23069
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 6730 23100 6736 23112
rect 6691 23072 6736 23100
rect 6730 23060 6736 23072
rect 6788 23060 6794 23112
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23100 19487 23103
rect 19610 23100 19616 23112
rect 19475 23072 19616 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 19610 23060 19616 23072
rect 19668 23100 19674 23112
rect 19886 23100 19892 23112
rect 19668 23072 19892 23100
rect 19668 23060 19674 23072
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 20438 23100 20444 23112
rect 20399 23072 20444 23100
rect 20438 23060 20444 23072
rect 20496 23060 20502 23112
rect 21266 23100 21272 23112
rect 21227 23072 21272 23100
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23100 21971 23103
rect 22204 23100 22232 23276
rect 22278 23100 22284 23112
rect 21959 23072 22284 23100
rect 21959 23069 21971 23072
rect 21913 23063 21971 23069
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 4798 23032 4804 23044
rect 4356 23004 4804 23032
rect 4249 22995 4307 23001
rect 4798 22992 4804 23004
rect 4856 22992 4862 23044
rect 5442 23032 5448 23044
rect 5403 23004 5448 23032
rect 5442 22992 5448 23004
rect 5500 22992 5506 23044
rect 16666 23032 16672 23044
rect 16627 23004 16672 23032
rect 16666 22992 16672 23004
rect 16724 22992 16730 23044
rect 16885 23035 16943 23041
rect 16885 23001 16897 23035
rect 16931 23032 16943 23035
rect 17218 23032 17224 23044
rect 16931 23004 17224 23032
rect 16931 23001 16943 23004
rect 16885 22995 16943 23001
rect 17218 22992 17224 23004
rect 17276 23032 17282 23044
rect 17497 23035 17555 23041
rect 17276 23004 17448 23032
rect 17276 22992 17282 23004
rect 3142 22924 3148 22976
rect 3200 22964 3206 22976
rect 3973 22967 4031 22973
rect 3973 22964 3985 22967
rect 3200 22936 3985 22964
rect 3200 22924 3206 22936
rect 3973 22933 3985 22936
rect 4019 22933 4031 22967
rect 3973 22927 4031 22933
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 5077 22967 5135 22973
rect 5077 22964 5089 22967
rect 4672 22936 5089 22964
rect 4672 22924 4678 22936
rect 5077 22933 5089 22936
rect 5123 22933 5135 22967
rect 5077 22927 5135 22933
rect 5166 22924 5172 22976
rect 5224 22964 5230 22976
rect 6549 22967 6607 22973
rect 6549 22964 6561 22967
rect 5224 22936 6561 22964
rect 5224 22924 5230 22936
rect 6549 22933 6561 22936
rect 6595 22933 6607 22967
rect 17420 22964 17448 23004
rect 17497 23001 17509 23035
rect 17543 23032 17555 23035
rect 18322 23032 18328 23044
rect 17543 23004 18328 23032
rect 17543 23001 17555 23004
rect 17497 22995 17555 23001
rect 18322 22992 18328 23004
rect 18380 22992 18386 23044
rect 19058 22992 19064 23044
rect 19116 23032 19122 23044
rect 20898 23032 20904 23044
rect 19116 23004 20904 23032
rect 19116 22992 19122 23004
rect 20898 22992 20904 23004
rect 20956 22992 20962 23044
rect 17678 22964 17684 22976
rect 17420 22936 17684 22964
rect 6549 22927 6607 22933
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22964 18015 22967
rect 19518 22964 19524 22976
rect 18003 22936 19524 22964
rect 18003 22933 18015 22936
rect 17957 22927 18015 22933
rect 19518 22924 19524 22936
rect 19576 22924 19582 22976
rect 19794 22964 19800 22976
rect 19707 22936 19800 22964
rect 19794 22924 19800 22936
rect 19852 22964 19858 22976
rect 20717 22967 20775 22973
rect 20717 22964 20729 22967
rect 19852 22936 20729 22964
rect 19852 22924 19858 22936
rect 20717 22933 20729 22936
rect 20763 22964 20775 22967
rect 21266 22964 21272 22976
rect 20763 22936 21272 22964
rect 20763 22933 20775 22936
rect 20717 22927 20775 22933
rect 21266 22924 21272 22936
rect 21324 22924 21330 22976
rect 1104 22874 22976 22896
rect 1104 22822 6378 22874
rect 6430 22822 6442 22874
rect 6494 22822 6506 22874
rect 6558 22822 6570 22874
rect 6622 22822 6634 22874
rect 6686 22822 11806 22874
rect 11858 22822 11870 22874
rect 11922 22822 11934 22874
rect 11986 22822 11998 22874
rect 12050 22822 12062 22874
rect 12114 22822 17234 22874
rect 17286 22822 17298 22874
rect 17350 22822 17362 22874
rect 17414 22822 17426 22874
rect 17478 22822 17490 22874
rect 17542 22822 22662 22874
rect 22714 22822 22726 22874
rect 22778 22822 22790 22874
rect 22842 22822 22854 22874
rect 22906 22822 22918 22874
rect 22970 22822 22976 22874
rect 1104 22800 22976 22822
rect 5166 22760 5172 22772
rect 1863 22732 5172 22760
rect 1863 22701 1891 22732
rect 5166 22720 5172 22732
rect 5224 22720 5230 22772
rect 7098 22760 7104 22772
rect 7059 22732 7104 22760
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 18230 22760 18236 22772
rect 18191 22732 18236 22760
rect 18230 22720 18236 22732
rect 18288 22720 18294 22772
rect 18601 22763 18659 22769
rect 18601 22729 18613 22763
rect 18647 22760 18659 22763
rect 19288 22760 19294 22772
rect 18647 22732 19294 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 19288 22720 19294 22732
rect 19346 22720 19352 22772
rect 19702 22720 19708 22772
rect 19760 22760 19766 22772
rect 20070 22760 20076 22772
rect 19760 22732 19932 22760
rect 20031 22732 20076 22760
rect 19760 22720 19766 22732
rect 1848 22695 1906 22701
rect 1848 22661 1860 22695
rect 1894 22661 1906 22695
rect 1848 22655 1906 22661
rect 3418 22652 3424 22704
rect 3476 22692 3482 22704
rect 3789 22695 3847 22701
rect 3789 22692 3801 22695
rect 3476 22664 3801 22692
rect 3476 22652 3482 22664
rect 3789 22661 3801 22664
rect 3835 22692 3847 22695
rect 4433 22695 4491 22701
rect 4433 22692 4445 22695
rect 3835 22664 4445 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 4433 22661 4445 22664
rect 4479 22661 4491 22695
rect 4433 22655 4491 22661
rect 4649 22695 4707 22701
rect 4649 22661 4661 22695
rect 4695 22692 4707 22695
rect 6822 22692 6828 22704
rect 4695 22664 6828 22692
rect 4695 22661 4707 22664
rect 4649 22655 4707 22661
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 18248 22692 18276 22720
rect 19426 22692 19432 22704
rect 17696 22664 18276 22692
rect 18432 22664 19432 22692
rect 1578 22624 1584 22636
rect 1491 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22624 1642 22636
rect 2314 22624 2320 22636
rect 1636 22596 2320 22624
rect 1636 22584 1642 22596
rect 2314 22584 2320 22596
rect 2372 22584 2378 22636
rect 4062 22584 4068 22636
rect 4120 22624 4126 22636
rect 5905 22627 5963 22633
rect 5905 22624 5917 22627
rect 4120 22596 5917 22624
rect 4120 22584 4126 22596
rect 5905 22593 5917 22596
rect 5951 22624 5963 22627
rect 6086 22624 6092 22636
rect 5951 22596 6092 22624
rect 5951 22593 5963 22596
rect 5905 22587 5963 22593
rect 6086 22584 6092 22596
rect 6144 22584 6150 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 8110 22624 8116 22636
rect 6687 22596 8116 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 2682 22516 2688 22568
rect 2740 22556 2746 22568
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 2740 22528 3433 22556
rect 2740 22516 2746 22528
rect 3421 22525 3433 22528
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 6656 22556 6684 22587
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 17696 22633 17724 22664
rect 18432 22633 18460 22664
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22593 17555 22627
rect 17497 22587 17555 22593
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 5408 22528 6684 22556
rect 17512 22556 17540 22587
rect 17862 22556 17868 22568
rect 17512 22528 17868 22556
rect 5408 22516 5414 22528
rect 17862 22516 17868 22528
rect 17920 22556 17926 22568
rect 18156 22556 18184 22587
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 19242 22624 19248 22636
rect 18748 22596 19248 22624
rect 18748 22584 18754 22596
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 19352 22633 19380 22664
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 19904 22692 19932 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 20162 22720 20168 22772
rect 20220 22760 20226 22772
rect 21634 22760 21640 22772
rect 20220 22732 21640 22760
rect 20220 22720 20226 22732
rect 21634 22720 21640 22732
rect 21692 22720 21698 22772
rect 22097 22763 22155 22769
rect 22097 22760 22109 22763
rect 22020 22732 22109 22760
rect 20714 22692 20720 22704
rect 19904 22664 20720 22692
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 21208 22695 21266 22701
rect 21208 22661 21220 22695
rect 21254 22692 21266 22695
rect 21450 22692 21456 22704
rect 21254 22664 21456 22692
rect 21254 22661 21266 22664
rect 21208 22655 21266 22661
rect 21450 22652 21456 22664
rect 21508 22652 21514 22704
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22624 19395 22627
rect 19613 22627 19671 22633
rect 19383 22596 19417 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 20162 22624 20168 22636
rect 19659 22596 20168 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 21818 22624 21824 22636
rect 20364 22596 21824 22624
rect 17920 22528 18184 22556
rect 17920 22516 17926 22528
rect 2314 22380 2320 22432
rect 2372 22420 2378 22432
rect 2700 22420 2728 22516
rect 2866 22448 2872 22500
rect 2924 22488 2930 22500
rect 2961 22491 3019 22497
rect 2961 22488 2973 22491
rect 2924 22460 2973 22488
rect 2924 22448 2930 22460
rect 2961 22457 2973 22460
rect 3007 22457 3019 22491
rect 2961 22451 3019 22457
rect 3878 22448 3884 22500
rect 3936 22488 3942 22500
rect 5261 22491 5319 22497
rect 5261 22488 5273 22491
rect 3936 22460 5273 22488
rect 3936 22448 3942 22460
rect 5261 22457 5273 22460
rect 5307 22457 5319 22491
rect 6730 22488 6736 22500
rect 5261 22451 5319 22457
rect 5736 22460 6736 22488
rect 2372 22392 2728 22420
rect 2372 22380 2378 22392
rect 3050 22380 3056 22432
rect 3108 22420 3114 22432
rect 3789 22423 3847 22429
rect 3789 22420 3801 22423
rect 3108 22392 3801 22420
rect 3108 22380 3114 22392
rect 3789 22389 3801 22392
rect 3835 22389 3847 22423
rect 3789 22383 3847 22389
rect 3973 22423 4031 22429
rect 3973 22389 3985 22423
rect 4019 22420 4031 22423
rect 4154 22420 4160 22432
rect 4019 22392 4160 22420
rect 4019 22389 4031 22392
rect 3973 22383 4031 22389
rect 4154 22380 4160 22392
rect 4212 22380 4218 22432
rect 4614 22420 4620 22432
rect 4575 22392 4620 22420
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 4801 22423 4859 22429
rect 4801 22389 4813 22423
rect 4847 22420 4859 22423
rect 5736 22420 5764 22460
rect 6730 22448 6736 22460
rect 6788 22448 6794 22500
rect 18156 22488 18184 22528
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 20364 22556 20392 22596
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 19567 22528 20392 22556
rect 21453 22559 21511 22565
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 21453 22525 21465 22559
rect 21499 22556 21511 22559
rect 21542 22556 21548 22568
rect 21499 22528 21548 22556
rect 21499 22525 21511 22528
rect 21453 22519 21511 22525
rect 21542 22516 21548 22528
rect 21600 22556 21606 22568
rect 22020 22556 22048 22732
rect 22097 22729 22109 22732
rect 22143 22729 22155 22763
rect 22097 22723 22155 22729
rect 22094 22584 22100 22636
rect 22152 22624 22158 22636
rect 22281 22627 22339 22633
rect 22281 22624 22293 22627
rect 22152 22596 22293 22624
rect 22152 22584 22158 22596
rect 22281 22593 22293 22596
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 21600 22528 22048 22556
rect 21600 22516 21606 22528
rect 18156 22460 20208 22488
rect 17586 22420 17592 22432
rect 4847 22392 5764 22420
rect 17547 22392 17592 22420
rect 4847 22389 4859 22392
rect 4801 22383 4859 22389
rect 17586 22380 17592 22392
rect 17644 22380 17650 22432
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19061 22423 19119 22429
rect 19061 22420 19073 22423
rect 18932 22392 19073 22420
rect 18932 22380 18938 22392
rect 19061 22389 19073 22392
rect 19107 22389 19119 22423
rect 19061 22383 19119 22389
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 20070 22420 20076 22432
rect 19668 22392 20076 22420
rect 19668 22380 19674 22392
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20180 22420 20208 22460
rect 21910 22420 21916 22432
rect 20180 22392 21916 22420
rect 21910 22380 21916 22392
rect 21968 22380 21974 22432
rect 1104 22330 22816 22352
rect 1104 22278 3664 22330
rect 3716 22278 3728 22330
rect 3780 22278 3792 22330
rect 3844 22278 3856 22330
rect 3908 22278 3920 22330
rect 3972 22278 9092 22330
rect 9144 22278 9156 22330
rect 9208 22278 9220 22330
rect 9272 22278 9284 22330
rect 9336 22278 9348 22330
rect 9400 22278 14520 22330
rect 14572 22278 14584 22330
rect 14636 22278 14648 22330
rect 14700 22278 14712 22330
rect 14764 22278 14776 22330
rect 14828 22278 19948 22330
rect 20000 22278 20012 22330
rect 20064 22278 20076 22330
rect 20128 22278 20140 22330
rect 20192 22278 20204 22330
rect 20256 22278 22816 22330
rect 1104 22256 22816 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 3418 22216 3424 22228
rect 2280 22188 3424 22216
rect 2280 22176 2286 22188
rect 3418 22176 3424 22188
rect 3476 22216 3482 22228
rect 4157 22219 4215 22225
rect 4157 22216 4169 22219
rect 3476 22188 4169 22216
rect 3476 22176 3482 22188
rect 4157 22185 4169 22188
rect 4203 22216 4215 22219
rect 4614 22216 4620 22228
rect 4203 22188 4620 22216
rect 4203 22185 4215 22188
rect 4157 22179 4215 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 5445 22219 5503 22225
rect 5445 22216 5457 22219
rect 5408 22188 5457 22216
rect 5408 22176 5414 22188
rect 5445 22185 5457 22188
rect 5491 22185 5503 22219
rect 5445 22179 5503 22185
rect 20257 22219 20315 22225
rect 20257 22185 20269 22219
rect 20303 22216 20315 22219
rect 20806 22216 20812 22228
rect 20303 22188 20812 22216
rect 20303 22185 20315 22188
rect 20257 22179 20315 22185
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 4341 22151 4399 22157
rect 4341 22117 4353 22151
rect 4387 22148 4399 22151
rect 4982 22148 4988 22160
rect 4387 22120 4988 22148
rect 4387 22117 4399 22120
rect 4341 22111 4399 22117
rect 4982 22108 4988 22120
rect 5040 22108 5046 22160
rect 16850 22108 16856 22160
rect 16908 22148 16914 22160
rect 19334 22148 19340 22160
rect 16908 22120 19340 22148
rect 16908 22108 16914 22120
rect 19334 22108 19340 22120
rect 19392 22108 19398 22160
rect 21082 22148 21088 22160
rect 19996 22120 21088 22148
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 4062 22040 4068 22092
rect 4120 22080 4126 22092
rect 4246 22080 4252 22092
rect 4120 22052 4252 22080
rect 4120 22040 4126 22052
rect 4246 22040 4252 22052
rect 4304 22040 4310 22092
rect 4706 22040 4712 22092
rect 4764 22080 4770 22092
rect 4893 22083 4951 22089
rect 4893 22080 4905 22083
rect 4764 22052 4905 22080
rect 4764 22040 4770 22052
rect 4893 22049 4905 22052
rect 4939 22049 4951 22083
rect 4893 22043 4951 22049
rect 6089 22083 6147 22089
rect 6089 22049 6101 22083
rect 6135 22080 6147 22083
rect 7282 22080 7288 22092
rect 6135 22052 7288 22080
rect 6135 22049 6147 22052
rect 6089 22043 6147 22049
rect 7282 22040 7288 22052
rect 7340 22040 7346 22092
rect 10594 22080 10600 22092
rect 10555 22052 10600 22080
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 18417 22083 18475 22089
rect 18417 22049 18429 22083
rect 18463 22080 18475 22083
rect 19996 22080 20024 22120
rect 21082 22108 21088 22120
rect 21140 22108 21146 22160
rect 21266 22080 21272 22092
rect 18463 22052 20024 22080
rect 21100 22052 21272 22080
rect 18463 22049 18475 22052
rect 18417 22043 18475 22049
rect 1854 22021 1860 22024
rect 1848 21975 1860 22021
rect 1912 22012 1918 22024
rect 1912 21984 1948 22012
rect 1854 21972 1860 21975
rect 1912 21972 1918 21984
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 3878 22012 3884 22024
rect 2464 21984 3884 22012
rect 2464 21972 2470 21984
rect 3878 21972 3884 21984
rect 3936 22012 3942 22024
rect 4798 22012 4804 22024
rect 3936 21984 4108 22012
rect 4759 21984 4804 22012
rect 3936 21972 3942 21984
rect 2866 21904 2872 21956
rect 2924 21944 2930 21956
rect 3973 21947 4031 21953
rect 3973 21944 3985 21947
rect 2924 21916 3985 21944
rect 2924 21904 2930 21916
rect 3973 21913 3985 21916
rect 4019 21913 4031 21947
rect 4080 21944 4108 21984
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 5684 21984 6561 22012
rect 5684 21972 5690 21984
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 22012 10747 22015
rect 11698 22012 11704 22024
rect 10735 21984 11704 22012
rect 10735 21981 10747 21984
rect 10689 21975 10747 21981
rect 11698 21972 11704 21984
rect 11756 21972 11762 22024
rect 18598 22012 18604 22024
rect 18559 21984 18604 22012
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18874 22012 18880 22024
rect 18835 21984 18880 22012
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19334 22012 19340 22024
rect 19260 21984 19340 22012
rect 4173 21947 4231 21953
rect 4173 21944 4185 21947
rect 4080 21916 4185 21944
rect 3973 21907 4031 21913
rect 4173 21913 4185 21916
rect 4219 21913 4231 21947
rect 4173 21907 4231 21913
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 19260 21944 19288 21984
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19886 22012 19892 22024
rect 19847 21984 19892 22012
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 21100 22012 21128 22052
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 20272 21984 21128 22012
rect 19978 21944 19984 21956
rect 17736 21916 19984 21944
rect 17736 21904 17742 21916
rect 19978 21904 19984 21916
rect 20036 21904 20042 21956
rect 20272 21888 20300 21984
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 22014 22015 22072 22021
rect 22014 22012 22026 22015
rect 21232 21984 22026 22012
rect 21232 21972 21238 21984
rect 22014 21981 22026 21984
rect 22060 21981 22072 22015
rect 22014 21975 22072 21981
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 20714 21944 20720 21956
rect 20456 21916 20720 21944
rect 2498 21836 2504 21888
rect 2556 21876 2562 21888
rect 2961 21879 3019 21885
rect 2961 21876 2973 21879
rect 2556 21848 2973 21876
rect 2556 21836 2562 21848
rect 2961 21845 2973 21848
rect 3007 21845 3019 21879
rect 2961 21839 3019 21845
rect 10321 21879 10379 21885
rect 10321 21845 10333 21879
rect 10367 21876 10379 21879
rect 10410 21876 10416 21888
rect 10367 21848 10416 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 10410 21836 10416 21848
rect 10468 21836 10474 21888
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17828 21848 17969 21876
rect 17828 21836 17834 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 18782 21876 18788 21888
rect 18743 21848 18788 21876
rect 17957 21839 18015 21845
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 20254 21876 20260 21888
rect 20215 21848 20260 21876
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 20456 21885 20484 21916
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 21542 21904 21548 21956
rect 21600 21944 21606 21956
rect 22296 21944 22324 21975
rect 21600 21916 22324 21944
rect 21600 21904 21606 21916
rect 20441 21879 20499 21885
rect 20441 21845 20453 21879
rect 20487 21845 20499 21879
rect 20441 21839 20499 21845
rect 20530 21836 20536 21888
rect 20588 21876 20594 21888
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20588 21848 20913 21876
rect 20588 21836 20594 21848
rect 20901 21845 20913 21848
rect 20947 21876 20959 21879
rect 21082 21876 21088 21888
rect 20947 21848 21088 21876
rect 20947 21845 20959 21848
rect 20901 21839 20959 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 2130 21672 2136 21684
rect 2091 21644 2136 21672
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 2590 21672 2596 21684
rect 2551 21644 2596 21672
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 2961 21675 3019 21681
rect 2961 21641 2973 21675
rect 3007 21672 3019 21675
rect 3142 21672 3148 21684
rect 3007 21644 3148 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 3142 21632 3148 21644
rect 3200 21632 3206 21684
rect 4341 21675 4399 21681
rect 4341 21641 4353 21675
rect 4387 21672 4399 21675
rect 4430 21672 4436 21684
rect 4387 21644 4436 21672
rect 4387 21641 4399 21644
rect 4341 21635 4399 21641
rect 4430 21632 4436 21644
rect 4488 21632 4494 21684
rect 4890 21672 4896 21684
rect 4803 21644 4896 21672
rect 4890 21632 4896 21644
rect 4948 21672 4954 21684
rect 5350 21672 5356 21684
rect 4948 21644 5356 21672
rect 4948 21632 4954 21644
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 18782 21632 18788 21684
rect 18840 21672 18846 21684
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 18840 21644 20821 21672
rect 18840 21632 18846 21644
rect 20809 21641 20821 21644
rect 20855 21641 20867 21675
rect 21266 21672 21272 21684
rect 20809 21635 20867 21641
rect 20916 21644 21272 21672
rect 1949 21607 2007 21613
rect 1949 21573 1961 21607
rect 1995 21604 2007 21607
rect 2222 21604 2228 21616
rect 1995 21576 2228 21604
rect 1995 21573 2007 21576
rect 1949 21567 2007 21573
rect 2222 21564 2228 21576
rect 2280 21564 2286 21616
rect 19426 21564 19432 21616
rect 19484 21604 19490 21616
rect 20254 21604 20260 21616
rect 19484 21576 20260 21604
rect 19484 21564 19490 21576
rect 20254 21564 20260 21576
rect 20312 21604 20318 21616
rect 20530 21604 20536 21616
rect 20312 21576 20536 21604
rect 20312 21564 20318 21576
rect 20530 21564 20536 21576
rect 20588 21564 20594 21616
rect 20714 21564 20720 21616
rect 20772 21604 20778 21616
rect 20916 21604 20944 21644
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 21082 21604 21088 21616
rect 20772 21576 20944 21604
rect 21043 21576 21088 21604
rect 20772 21564 20778 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 21177 21607 21235 21613
rect 21177 21573 21189 21607
rect 21223 21604 21235 21607
rect 22186 21604 22192 21616
rect 21223 21576 22192 21604
rect 21223 21573 21235 21576
rect 21177 21567 21235 21573
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 1581 21539 1639 21545
rect 1581 21505 1593 21539
rect 1627 21536 1639 21539
rect 2406 21536 2412 21548
rect 1627 21508 2412 21536
rect 1627 21505 1639 21508
rect 1581 21499 1639 21505
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 2774 21496 2780 21548
rect 2832 21536 2838 21548
rect 3053 21539 3111 21545
rect 2832 21508 2877 21536
rect 2832 21496 2838 21508
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 4154 21536 4160 21548
rect 4115 21508 4160 21536
rect 3053 21499 3111 21505
rect 2130 21428 2136 21480
rect 2188 21468 2194 21480
rect 3068 21468 3096 21499
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 9916 21508 9965 21536
rect 9916 21496 9922 21508
rect 9953 21505 9965 21508
rect 9999 21536 10011 21539
rect 10594 21536 10600 21548
rect 9999 21508 10600 21536
rect 9999 21505 10011 21508
rect 9953 21499 10011 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20806 21536 20812 21548
rect 19935 21508 20812 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20806 21496 20812 21508
rect 20864 21496 20870 21548
rect 20988 21539 21046 21545
rect 20988 21505 21000 21539
rect 21034 21505 21046 21539
rect 20988 21499 21046 21505
rect 2188 21440 3096 21468
rect 2188 21428 2194 21440
rect 3142 21428 3148 21480
rect 3200 21468 3206 21480
rect 3513 21471 3571 21477
rect 3513 21468 3525 21471
rect 3200 21440 3525 21468
rect 3200 21428 3206 21440
rect 3513 21437 3525 21440
rect 3559 21437 3571 21471
rect 19426 21468 19432 21480
rect 19387 21440 19432 21468
rect 3513 21431 3571 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 19978 21468 19984 21480
rect 19576 21440 19984 21468
rect 19576 21428 19582 21440
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21468 20407 21471
rect 20714 21468 20720 21480
rect 20395 21440 20720 21468
rect 20395 21437 20407 21440
rect 20349 21431 20407 21437
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 5810 21400 5816 21412
rect 1964 21372 5816 21400
rect 1964 21341 1992 21372
rect 5810 21360 5816 21372
rect 5868 21360 5874 21412
rect 19610 21360 19616 21412
rect 19668 21400 19674 21412
rect 20165 21403 20223 21409
rect 20165 21400 20177 21403
rect 19668 21372 20177 21400
rect 19668 21360 19674 21372
rect 20165 21369 20177 21372
rect 20211 21369 20223 21403
rect 20165 21363 20223 21369
rect 1949 21335 2007 21341
rect 1949 21301 1961 21335
rect 1995 21301 2007 21335
rect 1949 21295 2007 21301
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 10505 21335 10563 21341
rect 10505 21332 10517 21335
rect 10376 21304 10517 21332
rect 10376 21292 10382 21304
rect 10505 21301 10517 21304
rect 10551 21301 10563 21335
rect 10505 21295 10563 21301
rect 17770 21292 17776 21344
rect 17828 21332 17834 21344
rect 18693 21335 18751 21341
rect 18693 21332 18705 21335
rect 17828 21304 18705 21332
rect 17828 21292 17834 21304
rect 18693 21301 18705 21304
rect 18739 21301 18751 21335
rect 18693 21295 18751 21301
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 21008 21332 21036 21499
rect 21266 21496 21272 21548
rect 21324 21545 21330 21548
rect 21324 21539 21363 21545
rect 21351 21505 21363 21539
rect 21324 21499 21363 21505
rect 21324 21496 21330 21499
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 21508 21508 21553 21536
rect 21508 21496 21514 21508
rect 19300 21304 21036 21332
rect 19300 21292 19306 21304
rect 22002 21292 22008 21344
rect 22060 21332 22066 21344
rect 22281 21335 22339 21341
rect 22281 21332 22293 21335
rect 22060 21304 22293 21332
rect 22060 21292 22066 21304
rect 22281 21301 22293 21304
rect 22327 21301 22339 21335
rect 22281 21295 22339 21301
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 2130 21128 2136 21140
rect 2091 21100 2136 21128
rect 2130 21088 2136 21100
rect 2188 21088 2194 21140
rect 2777 21131 2835 21137
rect 2777 21097 2789 21131
rect 2823 21128 2835 21131
rect 3234 21128 3240 21140
rect 2823 21100 3240 21128
rect 2823 21097 2835 21100
rect 2777 21091 2835 21097
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 4065 21131 4123 21137
rect 4065 21097 4077 21131
rect 4111 21128 4123 21131
rect 4617 21131 4675 21137
rect 4617 21128 4629 21131
rect 4111 21100 4629 21128
rect 4111 21097 4123 21100
rect 4065 21091 4123 21097
rect 4617 21097 4629 21100
rect 4663 21128 4675 21131
rect 4890 21128 4896 21140
rect 4663 21100 4896 21128
rect 4663 21097 4675 21100
rect 4617 21091 4675 21097
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 11698 21128 11704 21140
rect 11659 21100 11704 21128
rect 11698 21088 11704 21100
rect 11756 21088 11762 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 19576 21100 20085 21128
rect 19576 21088 19582 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 20073 21091 20131 21097
rect 20257 21131 20315 21137
rect 20257 21097 20269 21131
rect 20303 21128 20315 21131
rect 20622 21128 20628 21140
rect 20303 21100 20628 21128
rect 20303 21097 20315 21100
rect 20257 21091 20315 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 21542 21128 21548 21140
rect 20916 21100 21548 21128
rect 1762 21020 1768 21072
rect 1820 21060 1826 21072
rect 2593 21063 2651 21069
rect 2593 21060 2605 21063
rect 1820 21032 2605 21060
rect 1820 21020 1826 21032
rect 2593 21029 2605 21032
rect 2639 21029 2651 21063
rect 2593 21023 2651 21029
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20992 1731 20995
rect 3326 20992 3332 21004
rect 1719 20964 3332 20992
rect 1719 20961 1731 20964
rect 1673 20955 1731 20961
rect 3326 20952 3332 20964
rect 3384 20952 3390 21004
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 6641 20995 6699 21001
rect 6641 20992 6653 20995
rect 4672 20964 6653 20992
rect 4672 20952 4678 20964
rect 6641 20961 6653 20964
rect 6687 20961 6699 20995
rect 6641 20955 6699 20961
rect 7374 20952 7380 21004
rect 7432 20992 7438 21004
rect 10318 20992 10324 21004
rect 7432 20964 10324 20992
rect 7432 20952 7438 20964
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 17770 20952 17776 21004
rect 17828 20992 17834 21004
rect 20916 21001 20944 21100
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22278 21128 22284 21140
rect 22239 21100 22284 21128
rect 22278 21088 22284 21100
rect 22336 21088 22342 21140
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 17828 20964 20913 20992
rect 17828 20952 17834 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 1762 20924 1768 20936
rect 1627 20896 1768 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 1857 20927 1915 20933
rect 1857 20893 1869 20927
rect 1903 20893 1915 20927
rect 1857 20887 1915 20893
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 4154 20924 4160 20936
rect 1995 20896 4160 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 1872 20856 1900 20887
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 2866 20856 2872 20868
rect 1872 20828 2872 20856
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 2961 20859 3019 20865
rect 2961 20825 2973 20859
rect 3007 20856 3019 20859
rect 4632 20856 4660 20952
rect 6733 20927 6791 20933
rect 6733 20893 6745 20927
rect 6779 20924 6791 20927
rect 8754 20924 8760 20936
rect 6779 20896 8760 20924
rect 6779 20893 6791 20896
rect 6733 20887 6791 20893
rect 8754 20884 8760 20896
rect 8812 20884 8818 20936
rect 10410 20884 10416 20936
rect 10468 20924 10474 20936
rect 10577 20927 10635 20933
rect 10577 20924 10589 20927
rect 10468 20896 10589 20924
rect 10468 20884 10474 20896
rect 10577 20893 10589 20896
rect 10623 20893 10635 20927
rect 10577 20887 10635 20893
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 18923 20896 19441 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19429 20893 19441 20896
rect 19475 20924 19487 20927
rect 19702 20924 19708 20936
rect 19475 20896 19708 20924
rect 19475 20893 19487 20896
rect 19429 20887 19487 20893
rect 19702 20884 19708 20896
rect 19760 20884 19766 20936
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21157 20927 21215 20933
rect 21157 20924 21169 20927
rect 21048 20896 21169 20924
rect 21048 20884 21054 20896
rect 21157 20893 21169 20896
rect 21203 20893 21215 20927
rect 21157 20887 21215 20893
rect 3007 20828 4660 20856
rect 3007 20825 3019 20828
rect 2961 20819 3019 20825
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 20225 20859 20283 20865
rect 20225 20856 20237 20859
rect 19852 20828 20237 20856
rect 19852 20816 19858 20828
rect 20225 20825 20237 20828
rect 20271 20825 20283 20859
rect 20225 20819 20283 20825
rect 20441 20859 20499 20865
rect 20441 20825 20453 20859
rect 20487 20856 20499 20859
rect 21634 20856 21640 20868
rect 20487 20828 21640 20856
rect 20487 20825 20499 20828
rect 20441 20819 20499 20825
rect 21634 20816 21640 20828
rect 21692 20816 21698 20868
rect 2761 20791 2819 20797
rect 2761 20757 2773 20791
rect 2807 20788 2819 20791
rect 3418 20788 3424 20800
rect 2807 20760 3424 20788
rect 2807 20757 2819 20760
rect 2761 20751 2819 20757
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 7098 20788 7104 20800
rect 7059 20760 7104 20788
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 19610 20788 19616 20800
rect 18380 20760 19616 20788
rect 18380 20748 18386 20760
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 1581 20587 1639 20593
rect 1581 20553 1593 20587
rect 1627 20584 1639 20587
rect 1946 20584 1952 20596
rect 1627 20556 1952 20584
rect 1627 20553 1639 20556
rect 1581 20547 1639 20553
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 3237 20587 3295 20593
rect 3237 20553 3249 20587
rect 3283 20584 3295 20587
rect 4798 20584 4804 20596
rect 3283 20556 4804 20584
rect 3283 20553 3295 20556
rect 3237 20547 3295 20553
rect 4798 20544 4804 20556
rect 4856 20544 4862 20596
rect 14553 20587 14611 20593
rect 14553 20553 14565 20587
rect 14599 20553 14611 20587
rect 14553 20547 14611 20553
rect 1762 20516 1768 20528
rect 1723 20488 1768 20516
rect 1762 20476 1768 20488
rect 1820 20476 1826 20528
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 7622 20519 7680 20525
rect 7622 20516 7634 20519
rect 7156 20488 7634 20516
rect 7156 20476 7162 20488
rect 7622 20485 7634 20488
rect 7668 20485 7680 20519
rect 7622 20479 7680 20485
rect 13848 20519 13906 20525
rect 13848 20485 13860 20519
rect 13894 20516 13906 20519
rect 14568 20516 14596 20547
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21285 20587 21343 20593
rect 21285 20584 21297 20587
rect 20956 20556 21297 20584
rect 20956 20544 20962 20556
rect 21285 20553 21297 20556
rect 21331 20553 21343 20587
rect 21285 20547 21343 20553
rect 21453 20587 21511 20593
rect 21453 20553 21465 20587
rect 21499 20584 21511 20587
rect 21726 20584 21732 20596
rect 21499 20556 21732 20584
rect 21499 20553 21511 20556
rect 21453 20547 21511 20553
rect 21726 20544 21732 20556
rect 21784 20544 21790 20596
rect 13894 20488 14596 20516
rect 13894 20485 13906 20488
rect 13848 20479 13906 20485
rect 20530 20476 20536 20528
rect 20588 20516 20594 20528
rect 21085 20519 21143 20525
rect 21085 20516 21097 20519
rect 20588 20488 21097 20516
rect 20588 20476 20594 20488
rect 21085 20485 21097 20488
rect 21131 20485 21143 20519
rect 21085 20479 21143 20485
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2314 20448 2320 20460
rect 1995 20420 2320 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2314 20408 2320 20420
rect 2372 20408 2378 20460
rect 3050 20448 3056 20460
rect 3011 20420 3056 20448
rect 3050 20408 3056 20420
rect 3108 20448 3114 20460
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3108 20420 3709 20448
rect 3108 20408 3114 20420
rect 3697 20417 3709 20420
rect 3743 20417 3755 20451
rect 7374 20448 7380 20460
rect 7335 20420 7380 20448
rect 3697 20411 3755 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 13354 20448 13360 20460
rect 12728 20420 13360 20448
rect 10594 20272 10600 20324
rect 10652 20312 10658 20324
rect 12728 20321 12756 20420
rect 13354 20408 13360 20420
rect 13412 20448 13418 20460
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 13412 20420 14933 20448
rect 13412 20408 13418 20420
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20346 20448 20352 20460
rect 20027 20420 20352 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20496 20420 20637 20448
rect 20496 20408 20502 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 16850 20380 16856 20392
rect 15059 20352 16856 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 12713 20315 12771 20321
rect 10652 20284 12664 20312
rect 10652 20272 10658 20284
rect 2406 20244 2412 20256
rect 2367 20216 2412 20244
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 8754 20244 8760 20256
rect 8667 20216 8760 20244
rect 8754 20204 8760 20216
rect 8812 20244 8818 20256
rect 12526 20244 12532 20256
rect 8812 20216 12532 20244
rect 8812 20204 8818 20216
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 12636 20244 12664 20284
rect 12713 20281 12725 20315
rect 12759 20281 12771 20315
rect 12713 20275 12771 20281
rect 14108 20244 14136 20343
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 14274 20244 14280 20256
rect 12636 20216 14280 20244
rect 14274 20204 14280 20216
rect 14332 20244 14338 20256
rect 17770 20244 17776 20256
rect 14332 20216 17776 20244
rect 14332 20204 14338 20216
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 22278 20244 22284 20256
rect 22239 20216 22284 20244
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 14274 20040 14280 20052
rect 14235 20012 14280 20040
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 21177 20043 21235 20049
rect 21177 20040 21189 20043
rect 20864 20012 21189 20040
rect 20864 20000 20870 20012
rect 21177 20009 21189 20012
rect 21223 20009 21235 20043
rect 21910 20040 21916 20052
rect 21871 20012 21916 20040
rect 21177 20003 21235 20009
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 22244 20012 22293 20040
rect 22244 20000 22250 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 22281 20003 22339 20009
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19668 19876 21864 19904
rect 19668 19864 19674 19876
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 1581 19839 1639 19845
rect 1581 19836 1593 19839
rect 1544 19808 1593 19836
rect 1544 19796 1550 19808
rect 1581 19805 1593 19808
rect 1627 19805 1639 19839
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 1581 19799 1639 19805
rect 1596 19768 1624 19799
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19836 20775 19839
rect 21358 19836 21364 19848
rect 20763 19808 21364 19836
rect 20763 19805 20775 19808
rect 20717 19799 20775 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 21836 19845 21864 19876
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 2869 19771 2927 19777
rect 2869 19768 2881 19771
rect 1596 19740 2881 19768
rect 2869 19737 2881 19740
rect 2915 19737 2927 19771
rect 2869 19731 2927 19737
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 3418 19700 3424 19712
rect 1811 19672 3424 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 1854 19456 1860 19508
rect 1912 19496 1918 19508
rect 2225 19499 2283 19505
rect 2225 19496 2237 19499
rect 1912 19468 2237 19496
rect 1912 19456 1918 19468
rect 2225 19465 2237 19468
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 11756 19468 13584 19496
rect 11756 19456 11762 19468
rect 2406 19360 2412 19372
rect 2367 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19320 2470 19372
rect 12388 19369 12394 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11195 19332 11713 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 12345 19363 12394 19369
rect 12345 19329 12357 19363
rect 12391 19329 12394 19363
rect 12345 19323 12394 19329
rect 12388 19320 12394 19323
rect 12446 19320 12452 19372
rect 12526 19369 12532 19372
rect 12504 19363 12532 19369
rect 12504 19329 12516 19363
rect 12504 19323 12532 19329
rect 12526 19320 12532 19323
rect 12584 19320 12590 19372
rect 13354 19360 13360 19372
rect 13315 19332 13360 19360
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 13556 19369 13584 19468
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22002 19360 22008 19372
rect 21499 19332 22008 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22002 19320 22008 19332
rect 22060 19360 22066 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 22060 19332 22293 19360
rect 22060 19320 22066 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22281 19323 22339 19329
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 12621 19295 12679 19301
rect 12621 19292 12633 19295
rect 9548 19264 12633 19292
rect 9548 19252 9554 19264
rect 12621 19261 12633 19264
rect 12667 19261 12679 19295
rect 12621 19255 12679 19261
rect 12820 19264 17632 19292
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2774 19116 2780 19168
rect 2832 19156 2838 19168
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 2832 19128 2881 19156
rect 2832 19116 2838 19128
rect 2869 19125 2881 19128
rect 2915 19125 2927 19159
rect 10962 19156 10968 19168
rect 10923 19128 10968 19156
rect 2869 19119 2927 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 12820 19156 12848 19264
rect 12897 19227 12955 19233
rect 12897 19193 12909 19227
rect 12943 19224 12955 19227
rect 17604 19224 17632 19264
rect 22097 19227 22155 19233
rect 22097 19224 22109 19227
rect 12943 19196 17540 19224
rect 17604 19196 22109 19224
rect 12943 19193 12955 19196
rect 12897 19187 12955 19193
rect 12308 19128 12848 19156
rect 17512 19156 17540 19196
rect 22097 19193 22109 19196
rect 22143 19193 22155 19227
rect 22097 19187 22155 19193
rect 22186 19156 22192 19168
rect 17512 19128 22192 19156
rect 12308 19116 12314 19128
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18952 2007 18955
rect 3050 18952 3056 18964
rect 1995 18924 3056 18952
rect 1995 18921 2007 18924
rect 1949 18915 2007 18921
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 21542 18952 21548 18964
rect 21503 18924 21548 18952
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 2685 18887 2743 18893
rect 2685 18884 2697 18887
rect 2056 18856 2697 18884
rect 2056 18757 2084 18856
rect 2685 18853 2697 18856
rect 2731 18884 2743 18887
rect 5718 18884 5724 18896
rect 2731 18856 5724 18884
rect 2731 18853 2743 18856
rect 2685 18847 2743 18853
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 6917 18819 6975 18825
rect 6917 18816 6929 18819
rect 6788 18788 6929 18816
rect 6788 18776 6794 18788
rect 6917 18785 6929 18788
rect 6963 18785 6975 18819
rect 6917 18779 6975 18785
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18748 2559 18751
rect 2774 18748 2780 18760
rect 2547 18720 2780 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 3326 18748 3332 18760
rect 3287 18720 3332 18748
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18748 7067 18751
rect 9490 18748 9496 18760
rect 7055 18720 9496 18748
rect 7055 18717 7067 18720
rect 7009 18711 7067 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 22278 18748 22284 18760
rect 22239 18720 22284 18748
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 4614 18680 4620 18692
rect 1596 18652 4620 18680
rect 1596 18621 1624 18652
rect 4614 18640 4620 18652
rect 4672 18640 4678 18692
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 2866 18572 2872 18624
rect 2924 18612 2930 18624
rect 3145 18615 3203 18621
rect 3145 18612 3157 18615
rect 2924 18584 3157 18612
rect 2924 18572 2930 18584
rect 3145 18581 3157 18584
rect 3191 18581 3203 18615
rect 7374 18612 7380 18624
rect 7335 18584 7380 18612
rect 3145 18575 3203 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 3326 18408 3332 18420
rect 2179 18380 3332 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 9490 18408 9496 18420
rect 9263 18380 9496 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 1949 18343 2007 18349
rect 1949 18309 1961 18343
rect 1995 18340 2007 18343
rect 2222 18340 2228 18352
rect 1995 18312 2228 18340
rect 1995 18309 2007 18312
rect 1949 18303 2007 18309
rect 2222 18300 2228 18312
rect 2280 18300 2286 18352
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 8082 18343 8140 18349
rect 8082 18340 8094 18343
rect 7432 18312 8094 18340
rect 7432 18300 7438 18312
rect 8082 18309 8094 18312
rect 8128 18309 8140 18343
rect 8082 18303 8140 18309
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 2958 18272 2964 18284
rect 2919 18244 2964 18272
rect 2777 18235 2835 18241
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18204 1639 18207
rect 2314 18204 2320 18216
rect 1627 18176 2320 18204
rect 1627 18173 1639 18176
rect 1581 18167 1639 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2792 18204 2820 18235
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 3108 18244 3153 18272
rect 3108 18232 3114 18244
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7524 18244 7849 18272
rect 7524 18232 7530 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 3326 18204 3332 18216
rect 2792 18176 3332 18204
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 2038 18096 2044 18148
rect 2096 18136 2102 18148
rect 2593 18139 2651 18145
rect 2593 18136 2605 18139
rect 2096 18108 2605 18136
rect 2096 18096 2102 18108
rect 2593 18105 2605 18108
rect 2639 18105 2651 18139
rect 22278 18136 22284 18148
rect 22239 18108 22284 18136
rect 2593 18099 2651 18105
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17864 22155 17867
rect 22186 17864 22192 17876
rect 22143 17836 22192 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 22186 17824 22192 17836
rect 22244 17824 22250 17876
rect 1486 17620 1492 17672
rect 1544 17660 1550 17672
rect 1581 17663 1639 17669
rect 1581 17660 1593 17663
rect 1544 17632 1593 17660
rect 1544 17620 1550 17632
rect 1581 17629 1593 17632
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 2648 17632 4169 17660
rect 2648 17620 2654 17632
rect 4157 17629 4169 17632
rect 4203 17629 4215 17663
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4157 17623 4215 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17660 21695 17663
rect 22278 17660 22284 17672
rect 21683 17632 22284 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 1826 17595 1884 17601
rect 1826 17592 1838 17595
rect 1728 17564 1838 17592
rect 1728 17552 1734 17564
rect 1826 17561 1838 17564
rect 1872 17561 1884 17595
rect 1826 17555 1884 17561
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 3973 17595 4031 17601
rect 3973 17592 3985 17595
rect 3292 17564 3985 17592
rect 3292 17552 3298 17564
rect 3973 17561 3985 17564
rect 4019 17592 4031 17595
rect 5810 17592 5816 17604
rect 4019 17564 5816 17592
rect 4019 17561 4031 17564
rect 3973 17555 4031 17561
rect 5810 17552 5816 17564
rect 5868 17552 5874 17604
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 2961 17527 3019 17533
rect 2961 17524 2973 17527
rect 2740 17496 2973 17524
rect 2740 17484 2746 17496
rect 2961 17493 2973 17496
rect 3007 17493 3019 17527
rect 4338 17524 4344 17536
rect 4299 17496 4344 17524
rect 2961 17487 3019 17493
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 4801 17527 4859 17533
rect 4801 17524 4813 17527
rect 4488 17496 4813 17524
rect 4488 17484 4494 17496
rect 4801 17493 4813 17496
rect 4847 17493 4859 17527
rect 4801 17487 4859 17493
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 2958 17280 2964 17292
rect 3016 17320 3022 17332
rect 5166 17320 5172 17332
rect 3016 17292 5172 17320
rect 3016 17280 3022 17292
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 1848 17255 1906 17261
rect 1848 17221 1860 17255
rect 1894 17252 1906 17255
rect 4430 17252 4436 17264
rect 1894 17224 4436 17252
rect 1894 17221 1906 17224
rect 1848 17215 1906 17221
rect 4430 17212 4436 17224
rect 4488 17212 4494 17264
rect 3418 17184 3424 17196
rect 3379 17156 3424 17184
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 3568 17156 4537 17184
rect 3568 17144 3574 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4525 17147 4583 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 3142 17076 3148 17128
rect 3200 17116 3206 17128
rect 4816 17116 4844 17147
rect 3200 17088 4844 17116
rect 3200 17076 3206 17088
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 3016 17020 3709 17048
rect 3016 17008 3022 17020
rect 3697 17017 3709 17020
rect 3743 17017 3755 17051
rect 3697 17011 3755 17017
rect 4154 17008 4160 17060
rect 4212 17048 4218 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 4212 17020 5273 17048
rect 4212 17008 4218 17020
rect 5261 17017 5273 17020
rect 5307 17017 5319 17051
rect 22278 17048 22284 17060
rect 22239 17020 22284 17048
rect 5261 17011 5319 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 4062 16980 4068 16992
rect 3927 16952 4068 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 4304 16952 4353 16980
rect 4304 16940 4310 16952
rect 4341 16949 4353 16952
rect 4387 16949 4399 16983
rect 4341 16943 4399 16949
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 7466 16980 7472 16992
rect 4948 16952 7472 16980
rect 4948 16940 4954 16952
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 1578 16776 1584 16788
rect 1491 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16776 1642 16788
rect 2958 16776 2964 16788
rect 1636 16748 2964 16776
rect 1636 16736 1642 16748
rect 2958 16736 2964 16748
rect 3016 16776 3022 16788
rect 4338 16776 4344 16788
rect 3016 16748 4108 16776
rect 4299 16748 4344 16776
rect 3016 16736 3022 16748
rect 1596 16649 1624 16736
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 3973 16643 4031 16649
rect 3973 16640 3985 16643
rect 3476 16612 3985 16640
rect 3476 16600 3482 16612
rect 3973 16609 3985 16612
rect 4019 16609 4031 16643
rect 4080 16640 4108 16748
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5994 16776 6000 16788
rect 5955 16748 6000 16776
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 4525 16711 4583 16717
rect 4525 16677 4537 16711
rect 4571 16708 4583 16711
rect 6086 16708 6092 16720
rect 4571 16680 6092 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 4890 16640 4896 16652
rect 4080 16612 4896 16640
rect 3973 16603 4031 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 6012 16612 6868 16640
rect 6012 16584 6040 16612
rect 1854 16581 1860 16584
rect 1848 16535 1860 16581
rect 1912 16572 1918 16584
rect 1912 16544 1948 16572
rect 1854 16532 1860 16535
rect 1912 16532 1918 16544
rect 2222 16532 2228 16584
rect 2280 16572 2286 16584
rect 4338 16572 4344 16584
rect 2280 16544 4344 16572
rect 2280 16532 2286 16544
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 5534 16572 5540 16584
rect 5000 16544 5540 16572
rect 5000 16513 5028 16544
rect 5534 16532 5540 16544
rect 5592 16572 5598 16584
rect 5994 16572 6000 16584
rect 5592 16544 6000 16572
rect 5592 16532 5598 16544
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6840 16581 6868 16612
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 22060 16612 22293 16640
rect 22060 16600 22066 16612
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 22281 16603 22339 16609
rect 6641 16575 6699 16581
rect 6641 16572 6653 16575
rect 6196 16544 6653 16572
rect 4985 16507 5043 16513
rect 4985 16504 4997 16507
rect 3068 16476 4997 16504
rect 3068 16448 3096 16476
rect 4985 16473 4997 16476
rect 5031 16473 5043 16507
rect 5166 16504 5172 16516
rect 5127 16476 5172 16504
rect 4985 16467 5043 16473
rect 5166 16464 5172 16476
rect 5224 16504 5230 16516
rect 6196 16513 6224 16544
rect 6641 16541 6653 16544
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 6181 16507 6239 16513
rect 6181 16504 6193 16507
rect 5224 16476 6193 16504
rect 5224 16464 5230 16476
rect 6181 16473 6193 16476
rect 6227 16473 6239 16507
rect 6181 16467 6239 16473
rect 2961 16439 3019 16445
rect 2961 16405 2973 16439
rect 3007 16436 3019 16439
rect 3050 16436 3056 16448
rect 3007 16408 3056 16436
rect 3007 16405 3019 16408
rect 2961 16399 3019 16405
rect 3050 16396 3056 16408
rect 3108 16396 3114 16448
rect 4338 16436 4344 16448
rect 4251 16408 4344 16436
rect 4338 16396 4344 16408
rect 4396 16436 4402 16448
rect 4798 16436 4804 16448
rect 4396 16408 4804 16436
rect 4396 16396 4402 16408
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 5353 16439 5411 16445
rect 5353 16436 5365 16439
rect 5316 16408 5365 16436
rect 5316 16396 5322 16408
rect 5353 16405 5365 16408
rect 5399 16405 5411 16439
rect 5810 16436 5816 16448
rect 5771 16408 5816 16436
rect 5353 16399 5411 16405
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 5994 16445 6000 16448
rect 5981 16439 6000 16445
rect 5981 16405 5993 16439
rect 5981 16399 6000 16405
rect 5994 16396 6000 16399
rect 6052 16396 6058 16448
rect 6270 16396 6276 16448
rect 6328 16436 6334 16448
rect 6641 16439 6699 16445
rect 6641 16436 6653 16439
rect 6328 16408 6653 16436
rect 6328 16396 6334 16408
rect 6641 16405 6653 16408
rect 6687 16405 6699 16439
rect 6641 16399 6699 16405
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 1581 16235 1639 16241
rect 1581 16201 1593 16235
rect 1627 16232 1639 16235
rect 2590 16232 2596 16244
rect 1627 16204 2596 16232
rect 1627 16201 1639 16204
rect 1581 16195 1639 16201
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3384 16204 3433 16232
rect 3384 16192 3390 16204
rect 3421 16201 3433 16204
rect 3467 16232 3479 16235
rect 5994 16232 6000 16244
rect 3467 16204 6000 16232
rect 3467 16201 3479 16204
rect 3421 16195 3479 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 22281 16235 22339 16241
rect 22281 16232 22293 16235
rect 22152 16204 22293 16232
rect 22152 16192 22158 16204
rect 22281 16201 22293 16204
rect 22327 16201 22339 16235
rect 22281 16195 22339 16201
rect 2716 16167 2774 16173
rect 2716 16133 2728 16167
rect 2762 16164 2774 16167
rect 5902 16164 5908 16176
rect 2762 16136 5908 16164
rect 2762 16133 2774 16136
rect 2716 16127 2774 16133
rect 5902 16124 5908 16136
rect 5960 16124 5966 16176
rect 6178 16124 6184 16176
rect 6236 16164 6242 16176
rect 6701 16167 6759 16173
rect 6701 16164 6713 16167
rect 6236 16136 6713 16164
rect 6236 16124 6242 16136
rect 6701 16133 6713 16136
rect 6747 16133 6759 16167
rect 6914 16164 6920 16176
rect 6875 16136 6920 16164
rect 6701 16127 6759 16133
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 2958 16096 2964 16108
rect 2919 16068 2964 16096
rect 2958 16056 2964 16068
rect 3016 16056 3022 16108
rect 4545 16099 4603 16105
rect 4545 16065 4557 16099
rect 4591 16096 4603 16099
rect 6546 16096 6552 16108
rect 4591 16068 6552 16096
rect 4591 16065 4603 16068
rect 4545 16059 4603 16065
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 22094 16096 22100 16108
rect 21499 16068 22100 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 4890 16028 4896 16040
rect 4847 16000 4896 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 5534 16028 5540 16040
rect 5368 16000 5540 16028
rect 5368 15969 5396 16000
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 5718 16028 5724 16040
rect 5679 16000 5724 16028
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 5353 15963 5411 15969
rect 5353 15929 5365 15963
rect 5399 15929 5411 15963
rect 5353 15923 5411 15929
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 4212 15864 5273 15892
rect 4212 15852 4218 15864
rect 5261 15861 5273 15864
rect 5307 15861 5319 15895
rect 5261 15855 5319 15861
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 5592 15864 6561 15892
rect 5592 15852 5598 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6730 15892 6736 15904
rect 6691 15864 6736 15892
rect 6549 15855 6607 15861
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3234 15688 3240 15700
rect 2832 15660 3240 15688
rect 2832 15648 2838 15660
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 4617 15691 4675 15697
rect 4617 15657 4629 15691
rect 4663 15688 4675 15691
rect 4706 15688 4712 15700
rect 4663 15660 4712 15688
rect 4663 15657 4675 15660
rect 4617 15651 4675 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 5074 15688 5080 15700
rect 5035 15660 5080 15688
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 5902 15688 5908 15700
rect 5863 15660 5908 15688
rect 5902 15648 5908 15660
rect 5960 15648 5966 15700
rect 6546 15688 6552 15700
rect 6507 15660 6552 15688
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 4246 15620 4252 15632
rect 2746 15592 4252 15620
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 2746 15552 2774 15592
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 4798 15580 4804 15632
rect 4856 15620 4862 15632
rect 6730 15620 6736 15632
rect 4856 15592 6736 15620
rect 4856 15580 4862 15592
rect 2639 15524 2774 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 2958 15512 2964 15564
rect 3016 15552 3022 15564
rect 3234 15552 3240 15564
rect 3016 15524 3240 15552
rect 3016 15512 3022 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 4154 15552 4160 15564
rect 3988 15524 4160 15552
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 2406 15484 2412 15496
rect 2367 15456 2412 15484
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15453 2835 15487
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 2777 15447 2835 15453
rect 1762 15376 1768 15428
rect 1820 15416 1826 15428
rect 2792 15416 2820 15447
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3988 15493 4016 15524
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4614 15552 4620 15564
rect 4264 15524 4620 15552
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 4264 15493 4292 15524
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 6270 15552 6276 15564
rect 5276 15524 6276 15552
rect 4522 15493 4528 15496
rect 4249 15487 4307 15493
rect 4120 15456 4165 15484
rect 4120 15444 4126 15456
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 4479 15487 4528 15493
rect 4479 15453 4491 15487
rect 4525 15453 4528 15487
rect 4479 15447 4528 15453
rect 4522 15444 4528 15447
rect 4580 15444 4586 15496
rect 1820 15388 2820 15416
rect 1820 15376 1826 15388
rect 2958 15376 2964 15428
rect 3016 15416 3022 15428
rect 3326 15416 3332 15428
rect 3016 15388 3332 15416
rect 3016 15376 3022 15388
rect 3326 15376 3332 15388
rect 3384 15416 3390 15428
rect 5276 15425 5304 15524
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6086 15484 6092 15496
rect 6047 15456 6092 15484
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 4341 15419 4399 15425
rect 4341 15416 4353 15419
rect 3384 15388 4353 15416
rect 3384 15376 3390 15388
rect 4341 15385 4353 15388
rect 4387 15385 4399 15419
rect 4341 15379 4399 15385
rect 5245 15419 5304 15425
rect 5245 15385 5257 15419
rect 5291 15388 5304 15419
rect 5445 15419 5503 15425
rect 5291 15385 5303 15388
rect 5245 15379 5303 15385
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 6380 15416 6408 15592
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 10962 15484 10968 15496
rect 7699 15456 10968 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 22278 15484 22284 15496
rect 22239 15456 22284 15484
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 5491 15388 6408 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 1857 15351 1915 15357
rect 1857 15317 1869 15351
rect 1903 15348 1915 15351
rect 1946 15348 1952 15360
rect 1903 15320 1952 15348
rect 1903 15317 1915 15320
rect 1857 15311 1915 15317
rect 1946 15308 1952 15320
rect 2004 15348 2010 15360
rect 2222 15348 2228 15360
rect 2004 15320 2228 15348
rect 2004 15308 2010 15320
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 3602 15348 3608 15360
rect 2372 15320 3608 15348
rect 2372 15308 2378 15320
rect 3602 15308 3608 15320
rect 3660 15348 3666 15360
rect 6178 15348 6184 15360
rect 3660 15320 6184 15348
rect 3660 15308 3666 15320
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3973 15147 4031 15153
rect 3973 15144 3985 15147
rect 3568 15116 3985 15144
rect 3568 15104 3574 15116
rect 3973 15113 3985 15116
rect 4019 15113 4031 15147
rect 3973 15107 4031 15113
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 4982 15144 4988 15156
rect 4939 15116 4988 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15113 5411 15147
rect 5353 15107 5411 15113
rect 2590 15036 2596 15088
rect 2648 15036 2654 15088
rect 2716 15079 2774 15085
rect 2716 15045 2728 15079
rect 2762 15076 2774 15079
rect 5368 15076 5396 15107
rect 2762 15048 5396 15076
rect 2762 15045 2774 15048
rect 2716 15039 2774 15045
rect 2608 15008 2636 15036
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 2608 14980 3433 15008
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4062 15008 4068 15020
rect 3835 14980 4068 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 3326 14940 3332 14952
rect 3007 14912 3332 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 3326 14900 3332 14912
rect 3384 14940 3390 14952
rect 3510 14940 3516 14952
rect 3384 14912 3516 14940
rect 3384 14900 3390 14912
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 3620 14804 3648 14971
rect 3712 14940 3740 14971
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 15008 4491 15011
rect 5166 15008 5172 15020
rect 4479 14980 5172 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5534 15008 5540 15020
rect 5495 14980 5540 15008
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 4154 14940 4160 14952
rect 3712 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4798 14872 4804 14884
rect 4759 14844 4804 14872
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 22278 14872 22284 14884
rect 22239 14844 22284 14872
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 2648 14776 3648 14804
rect 2648 14764 2654 14776
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 4028 14572 4997 14600
rect 4028 14560 4034 14572
rect 4985 14569 4997 14572
rect 5031 14569 5043 14603
rect 4985 14563 5043 14569
rect 3234 14492 3240 14544
rect 3292 14532 3298 14544
rect 4801 14535 4859 14541
rect 4801 14532 4813 14535
rect 3292 14504 4813 14532
rect 3292 14492 3298 14504
rect 4801 14501 4813 14504
rect 4847 14501 4859 14535
rect 4801 14495 4859 14501
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3694 14464 3700 14476
rect 3007 14436 3700 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 4338 14464 4344 14476
rect 4299 14436 4344 14464
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 2705 14399 2763 14405
rect 2705 14365 2717 14399
rect 2751 14396 2763 14399
rect 2866 14396 2872 14408
rect 2751 14368 2872 14396
rect 2751 14365 2763 14368
rect 2705 14359 2763 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 3936 14368 5641 14396
rect 3936 14356 3942 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 3418 14288 3424 14340
rect 3476 14328 3482 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3476 14300 3985 14328
rect 3476 14288 3482 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4212 14300 4305 14328
rect 4212 14288 4218 14300
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 5169 14331 5227 14337
rect 5169 14328 5181 14331
rect 4856 14300 5181 14328
rect 4856 14288 4862 14300
rect 5169 14297 5181 14300
rect 5215 14297 5227 14331
rect 5169 14291 5227 14297
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 2682 14260 2688 14272
rect 1627 14232 2688 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 2682 14220 2688 14232
rect 2740 14260 2746 14272
rect 4172 14260 4200 14288
rect 2740 14232 4200 14260
rect 2740 14220 2746 14232
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 4959 14263 5017 14269
rect 4959 14260 4971 14263
rect 4672 14232 4971 14260
rect 4672 14220 4678 14232
rect 4959 14229 4971 14232
rect 5005 14229 5017 14263
rect 4959 14223 5017 14229
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 2958 14056 2964 14068
rect 2179 14028 2774 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 2746 13920 2774 14028
rect 2884 14028 2964 14056
rect 2884 13929 2912 14028
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4522 14056 4528 14068
rect 4483 14028 4528 14056
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 4540 13988 4568 14016
rect 2976 13960 4568 13988
rect 2976 13929 3004 13960
rect 2869 13923 2927 13929
rect 2746 13892 2820 13920
rect 2498 13812 2504 13864
rect 2556 13852 2562 13864
rect 2685 13855 2743 13861
rect 2685 13852 2697 13855
rect 2556 13824 2697 13852
rect 2556 13812 2562 13824
rect 2685 13821 2697 13824
rect 2731 13821 2743 13855
rect 2792 13852 2820 13892
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3384 13892 3617 13920
rect 3384 13880 3390 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 4246 13920 4252 13932
rect 3844 13892 4252 13920
rect 3844 13880 3850 13892
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4430 13920 4436 13932
rect 4391 13892 4436 13920
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 6730 13852 6736 13864
rect 2792 13824 6736 13852
rect 2685 13815 2743 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 22278 13852 22284 13864
rect 22239 13824 22284 13852
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13784 1639 13787
rect 2774 13784 2780 13796
rect 1627 13756 2780 13784
rect 1627 13753 1639 13756
rect 1581 13747 1639 13753
rect 2774 13744 2780 13756
rect 2832 13784 2838 13796
rect 3142 13784 3148 13796
rect 2832 13756 3148 13784
rect 2832 13744 2838 13756
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2038 13716 2044 13728
rect 1995 13688 2044 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 3786 13716 3792 13728
rect 2924 13688 3792 13716
rect 2924 13676 2930 13688
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1762 13512 1768 13524
rect 1719 13484 1768 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 2406 13512 2412 13524
rect 2179 13484 2412 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 2682 13512 2688 13524
rect 2516 13484 2688 13512
rect 2516 13376 2544 13484
rect 2682 13472 2688 13484
rect 2740 13512 2746 13524
rect 2777 13515 2835 13521
rect 2777 13512 2789 13515
rect 2740 13484 2789 13512
rect 2740 13472 2746 13484
rect 2777 13481 2789 13484
rect 2823 13481 2835 13515
rect 2777 13475 2835 13481
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 3326 13512 3332 13524
rect 3007 13484 3332 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 2866 13376 2872 13388
rect 1872 13348 2544 13376
rect 2700 13348 2872 13376
rect 1872 13317 1900 13348
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 1596 13240 1624 13271
rect 1946 13268 1952 13320
rect 2004 13308 2010 13320
rect 2700 13308 2728 13348
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 2004 13280 2049 13308
rect 2148 13280 2728 13308
rect 2004 13268 2010 13280
rect 2148 13240 2176 13280
rect 1596 13212 2176 13240
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2619 13243 2677 13249
rect 2619 13240 2631 13243
rect 2372 13212 2631 13240
rect 2372 13200 2378 13212
rect 2619 13209 2631 13212
rect 2665 13209 2677 13243
rect 3068 13240 3096 13484
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 4430 13512 4436 13524
rect 4203 13484 4436 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3568 13280 3985 13308
rect 3568 13268 3574 13280
rect 3973 13277 3985 13280
rect 4019 13308 4031 13311
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4019 13280 4629 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 22278 13308 22284 13320
rect 22239 13280 22284 13308
rect 4617 13271 4675 13277
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 2619 13203 2677 13209
rect 2746 13212 3096 13240
rect 2406 13132 2412 13184
rect 2464 13172 2470 13184
rect 2746 13172 2774 13212
rect 2464 13144 2774 13172
rect 2803 13175 2861 13181
rect 2464 13132 2470 13144
rect 2803 13141 2815 13175
rect 2849 13172 2861 13175
rect 3142 13172 3148 13184
rect 2849 13144 3148 13172
rect 2849 13141 2861 13144
rect 2803 13135 2861 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 2593 12971 2651 12977
rect 2593 12937 2605 12971
rect 2639 12968 2651 12971
rect 4614 12968 4620 12980
rect 2639 12940 4620 12968
rect 2639 12937 2651 12940
rect 2593 12931 2651 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 3142 12900 3148 12912
rect 1780 12872 3148 12900
rect 1780 12841 1808 12872
rect 3142 12860 3148 12872
rect 3200 12860 3206 12912
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 1765 12795 1823 12801
rect 1688 12696 1716 12795
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2866 12832 2872 12844
rect 2639 12804 2872 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3050 12832 3056 12844
rect 3011 12804 3056 12832
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3510 12792 3516 12844
rect 3568 12832 3574 12844
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3568 12804 3893 12832
rect 3568 12792 3574 12804
rect 3881 12801 3893 12804
rect 3927 12832 3939 12835
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 3927 12804 4353 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 3418 12764 3424 12776
rect 1995 12736 3424 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 2314 12696 2320 12708
rect 1688 12668 2320 12696
rect 2314 12656 2320 12668
rect 2372 12696 2378 12708
rect 2590 12696 2596 12708
rect 2372 12668 2596 12696
rect 2372 12656 2378 12668
rect 2590 12656 2596 12668
rect 2648 12656 2654 12708
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3200 12600 3709 12628
rect 3200 12588 3206 12600
rect 3697 12597 3709 12600
rect 3743 12597 3755 12631
rect 3697 12591 3755 12597
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1765 12427 1823 12433
rect 1765 12424 1777 12427
rect 1728 12396 1777 12424
rect 1728 12384 1734 12396
rect 1765 12393 1777 12396
rect 1811 12393 1823 12427
rect 1765 12387 1823 12393
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2774 12424 2780 12436
rect 2271 12396 2780 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 4062 12424 4068 12436
rect 3007 12396 4068 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 1946 12316 1952 12368
rect 2004 12356 2010 12368
rect 2976 12356 3004 12387
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 2004 12328 3004 12356
rect 2004 12316 2010 12328
rect 3234 12288 3240 12300
rect 1596 12260 3240 12288
rect 1596 12229 1624 12260
rect 3234 12248 3240 12260
rect 3292 12248 3298 12300
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2832 12192 2881 12220
rect 2832 12180 2838 12192
rect 2869 12189 2881 12192
rect 2915 12189 2927 12223
rect 22278 12220 22284 12232
rect 22239 12192 22284 12220
rect 2869 12183 2927 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 1673 11883 1731 11889
rect 1673 11849 1685 11883
rect 1719 11880 1731 11883
rect 2498 11880 2504 11892
rect 1719 11852 2504 11880
rect 1719 11849 1731 11852
rect 1673 11843 1731 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 3142 11812 3148 11824
rect 1780 11784 3148 11812
rect 1780 11753 1808 11784
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 1765 11707 1823 11713
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 22278 11608 22284 11620
rect 22239 11580 22284 11608
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1581 11135 1639 11141
rect 1581 11132 1593 11135
rect 1544 11104 1593 11132
rect 1544 11092 1550 11104
rect 1581 11101 1593 11104
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2774 10792 2780 10804
rect 1811 10764 2780 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10656 1642 10668
rect 2225 10659 2283 10665
rect 2225 10656 2237 10659
rect 1636 10628 2237 10656
rect 1636 10616 1642 10628
rect 2225 10625 2237 10628
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 22278 10520 22284 10532
rect 22239 10492 22284 10520
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 22278 10044 22284 10056
rect 22239 10016 22284 10044
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 1762 8956 1768 8968
rect 1723 8928 1768 8956
rect 1762 8916 1768 8928
rect 1820 8956 1826 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 1820 8928 2237 8956
rect 1820 8916 1826 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 22278 8956 22284 8968
rect 22239 8928 22284 8956
rect 2225 8919 2283 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 22278 8344 22284 8356
rect 22239 8316 22284 8344
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 22278 7256 22284 7268
rect 22239 7228 22284 7256
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 22278 6780 22284 6792
rect 22239 6752 22284 6780
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 7466 6304 7472 6316
rect 1903 6276 7472 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 22278 5692 22284 5704
rect 22239 5664 22284 5692
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 22278 5080 22284 5092
rect 22239 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 22278 3992 22284 4004
rect 22239 3964 22284 3992
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 22278 3516 22284 3528
rect 22239 3488 22284 3516
rect 22278 3476 22284 3488
rect 22336 3476 22342 3528
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 3976 27820 4028 27872
rect 7472 27820 7524 27872
rect 3664 27718 3716 27770
rect 3728 27718 3780 27770
rect 3792 27718 3844 27770
rect 3856 27718 3908 27770
rect 3920 27718 3972 27770
rect 9092 27718 9144 27770
rect 9156 27718 9208 27770
rect 9220 27718 9272 27770
rect 9284 27718 9336 27770
rect 9348 27718 9400 27770
rect 14520 27718 14572 27770
rect 14584 27718 14636 27770
rect 14648 27718 14700 27770
rect 14712 27718 14764 27770
rect 14776 27718 14828 27770
rect 19948 27718 20000 27770
rect 20012 27718 20064 27770
rect 20076 27718 20128 27770
rect 20140 27718 20192 27770
rect 20204 27718 20256 27770
rect 4068 27616 4120 27668
rect 7564 27616 7616 27668
rect 11980 27616 12032 27668
rect 6828 27548 6880 27600
rect 1768 27412 1820 27464
rect 3240 27480 3292 27532
rect 5264 27412 5316 27464
rect 5724 27412 5776 27464
rect 6092 27412 6144 27464
rect 6276 27344 6328 27396
rect 1860 27276 1912 27328
rect 2412 27319 2464 27328
rect 2412 27285 2421 27319
rect 2421 27285 2455 27319
rect 2455 27285 2464 27319
rect 2412 27276 2464 27285
rect 2964 27319 3016 27328
rect 2964 27285 2973 27319
rect 2973 27285 3007 27319
rect 3007 27285 3016 27319
rect 2964 27276 3016 27285
rect 4068 27319 4120 27328
rect 4068 27285 4077 27319
rect 4077 27285 4111 27319
rect 4111 27285 4120 27319
rect 4068 27276 4120 27285
rect 5356 27319 5408 27328
rect 5356 27285 5365 27319
rect 5365 27285 5399 27319
rect 5399 27285 5408 27319
rect 5356 27276 5408 27285
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 6828 27344 6880 27396
rect 6920 27344 6972 27396
rect 10324 27344 10376 27396
rect 10784 27344 10836 27396
rect 8392 27276 8444 27328
rect 10140 27276 10192 27328
rect 10692 27276 10744 27328
rect 11060 27344 11112 27396
rect 14464 27616 14516 27668
rect 14004 27548 14056 27600
rect 16948 27548 17000 27600
rect 19432 27548 19484 27600
rect 20352 27548 20404 27600
rect 12716 27523 12768 27532
rect 12716 27489 12725 27523
rect 12725 27489 12759 27523
rect 12759 27489 12768 27523
rect 12716 27480 12768 27489
rect 14188 27480 14240 27532
rect 12532 27455 12584 27464
rect 12532 27421 12541 27455
rect 12541 27421 12575 27455
rect 12575 27421 12584 27455
rect 12532 27412 12584 27421
rect 12900 27455 12952 27464
rect 12900 27421 12909 27455
rect 12909 27421 12943 27455
rect 12943 27421 12952 27455
rect 12900 27412 12952 27421
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 13268 27412 13320 27464
rect 14648 27480 14700 27532
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 17960 27412 18012 27464
rect 18604 27412 18656 27464
rect 20536 27412 20588 27464
rect 22100 27455 22152 27464
rect 22100 27421 22109 27455
rect 22109 27421 22143 27455
rect 22143 27421 22152 27455
rect 22100 27412 22152 27421
rect 13176 27344 13228 27396
rect 14648 27387 14700 27396
rect 11704 27276 11756 27328
rect 13452 27276 13504 27328
rect 14648 27353 14657 27387
rect 14657 27353 14691 27387
rect 14691 27353 14700 27387
rect 14648 27344 14700 27353
rect 15752 27344 15804 27396
rect 18144 27319 18196 27328
rect 18144 27285 18153 27319
rect 18153 27285 18187 27319
rect 18187 27285 18196 27319
rect 18144 27276 18196 27285
rect 21364 27319 21416 27328
rect 21364 27285 21373 27319
rect 21373 27285 21407 27319
rect 21407 27285 21416 27319
rect 21364 27276 21416 27285
rect 21824 27276 21876 27328
rect 6378 27174 6430 27226
rect 6442 27174 6494 27226
rect 6506 27174 6558 27226
rect 6570 27174 6622 27226
rect 6634 27174 6686 27226
rect 11806 27174 11858 27226
rect 11870 27174 11922 27226
rect 11934 27174 11986 27226
rect 11998 27174 12050 27226
rect 12062 27174 12114 27226
rect 17234 27174 17286 27226
rect 17298 27174 17350 27226
rect 17362 27174 17414 27226
rect 17426 27174 17478 27226
rect 17490 27174 17542 27226
rect 22662 27174 22714 27226
rect 22726 27174 22778 27226
rect 22790 27174 22842 27226
rect 22854 27174 22906 27226
rect 22918 27174 22970 27226
rect 5356 27072 5408 27124
rect 1584 27047 1636 27056
rect 1584 27013 1593 27047
rect 1593 27013 1627 27047
rect 1627 27013 1636 27047
rect 1584 27004 1636 27013
rect 3056 27004 3108 27056
rect 4068 27004 4120 27056
rect 2044 26936 2096 26988
rect 3516 26936 3568 26988
rect 4528 26979 4580 26988
rect 4528 26945 4537 26979
rect 4537 26945 4571 26979
rect 4571 26945 4580 26979
rect 4528 26936 4580 26945
rect 5172 26979 5224 26988
rect 5172 26945 5181 26979
rect 5181 26945 5215 26979
rect 5215 26945 5224 26979
rect 5172 26936 5224 26945
rect 7012 27004 7064 27056
rect 7656 27004 7708 27056
rect 7748 27004 7800 27056
rect 8024 27072 8076 27124
rect 9956 27072 10008 27124
rect 10048 27072 10100 27124
rect 11704 27072 11756 27124
rect 12532 27072 12584 27124
rect 14556 27115 14608 27124
rect 14556 27081 14565 27115
rect 14565 27081 14599 27115
rect 14599 27081 14608 27115
rect 14556 27072 14608 27081
rect 20536 27115 20588 27124
rect 20536 27081 20545 27115
rect 20545 27081 20579 27115
rect 20579 27081 20588 27115
rect 20536 27072 20588 27081
rect 8208 27004 8260 27056
rect 6828 26936 6880 26988
rect 11980 27004 12032 27056
rect 10876 26979 10928 26988
rect 5264 26868 5316 26920
rect 6644 26868 6696 26920
rect 10876 26945 10894 26979
rect 10894 26945 10928 26979
rect 10876 26936 10928 26945
rect 11520 26936 11572 26988
rect 13084 27004 13136 27056
rect 13176 26936 13228 26988
rect 13636 27004 13688 27056
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 18144 27004 18196 27056
rect 14004 26936 14056 26988
rect 16580 26936 16632 26988
rect 21916 27004 21968 27056
rect 20352 26979 20404 26988
rect 20352 26945 20361 26979
rect 20361 26945 20395 26979
rect 20395 26945 20404 26979
rect 20352 26936 20404 26945
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 8484 26800 8536 26852
rect 8944 26800 8996 26852
rect 1676 26732 1728 26784
rect 2504 26732 2556 26784
rect 2688 26732 2740 26784
rect 2872 26732 2924 26784
rect 5356 26775 5408 26784
rect 5356 26741 5365 26775
rect 5365 26741 5399 26775
rect 5399 26741 5408 26775
rect 5356 26732 5408 26741
rect 7012 26775 7064 26784
rect 7012 26741 7021 26775
rect 7021 26741 7055 26775
rect 7055 26741 7064 26775
rect 7012 26732 7064 26741
rect 7380 26732 7432 26784
rect 9496 26732 9548 26784
rect 11428 26868 11480 26920
rect 13084 26911 13136 26920
rect 13084 26877 13093 26911
rect 13093 26877 13127 26911
rect 13127 26877 13136 26911
rect 13084 26868 13136 26877
rect 11244 26732 11296 26784
rect 11612 26732 11664 26784
rect 14924 26800 14976 26852
rect 18144 26868 18196 26920
rect 20536 26868 20588 26920
rect 21088 26800 21140 26852
rect 12440 26732 12492 26784
rect 12900 26732 12952 26784
rect 13912 26732 13964 26784
rect 14648 26732 14700 26784
rect 17960 26775 18012 26784
rect 17960 26741 17969 26775
rect 17969 26741 18003 26775
rect 18003 26741 18012 26775
rect 17960 26732 18012 26741
rect 21456 26775 21508 26784
rect 21456 26741 21465 26775
rect 21465 26741 21499 26775
rect 21499 26741 21508 26775
rect 21456 26732 21508 26741
rect 21548 26732 21600 26784
rect 3664 26630 3716 26682
rect 3728 26630 3780 26682
rect 3792 26630 3844 26682
rect 3856 26630 3908 26682
rect 3920 26630 3972 26682
rect 9092 26630 9144 26682
rect 9156 26630 9208 26682
rect 9220 26630 9272 26682
rect 9284 26630 9336 26682
rect 9348 26630 9400 26682
rect 14520 26630 14572 26682
rect 14584 26630 14636 26682
rect 14648 26630 14700 26682
rect 14712 26630 14764 26682
rect 14776 26630 14828 26682
rect 19948 26630 20000 26682
rect 20012 26630 20064 26682
rect 20076 26630 20128 26682
rect 20140 26630 20192 26682
rect 20204 26630 20256 26682
rect 2044 26571 2096 26580
rect 2044 26537 2053 26571
rect 2053 26537 2087 26571
rect 2087 26537 2096 26571
rect 2044 26528 2096 26537
rect 4068 26528 4120 26580
rect 6736 26528 6788 26580
rect 6920 26571 6972 26580
rect 6920 26537 6929 26571
rect 6929 26537 6963 26571
rect 6963 26537 6972 26571
rect 6920 26528 6972 26537
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 7656 26528 7708 26580
rect 8208 26528 8260 26580
rect 2228 26460 2280 26512
rect 2780 26503 2832 26512
rect 2780 26469 2789 26503
rect 2789 26469 2823 26503
rect 2823 26469 2832 26503
rect 2780 26460 2832 26469
rect 7748 26460 7800 26512
rect 9680 26460 9732 26512
rect 9772 26460 9824 26512
rect 8668 26392 8720 26444
rect 10048 26571 10100 26580
rect 10048 26537 10057 26571
rect 10057 26537 10091 26571
rect 10091 26537 10100 26571
rect 10048 26528 10100 26537
rect 12808 26528 12860 26580
rect 14464 26571 14516 26580
rect 14464 26537 14473 26571
rect 14473 26537 14507 26571
rect 14507 26537 14516 26571
rect 14464 26528 14516 26537
rect 11980 26460 12032 26512
rect 12164 26460 12216 26512
rect 12348 26460 12400 26512
rect 13084 26460 13136 26512
rect 14280 26503 14332 26512
rect 14280 26469 14289 26503
rect 14289 26469 14323 26503
rect 14323 26469 14332 26503
rect 14280 26460 14332 26469
rect 14372 26460 14424 26512
rect 2412 26324 2464 26376
rect 5448 26367 5500 26376
rect 1584 26299 1636 26308
rect 1584 26265 1593 26299
rect 1593 26265 1627 26299
rect 1627 26265 1636 26299
rect 1584 26256 1636 26265
rect 2504 26256 2556 26308
rect 3240 26256 3292 26308
rect 3332 26256 3384 26308
rect 5448 26333 5457 26367
rect 5457 26333 5491 26367
rect 5491 26333 5500 26367
rect 5448 26324 5500 26333
rect 5724 26324 5776 26376
rect 6736 26367 6788 26376
rect 2964 26231 3016 26240
rect 2964 26197 2973 26231
rect 2973 26197 3007 26231
rect 3007 26197 3016 26231
rect 2964 26188 3016 26197
rect 3148 26188 3200 26240
rect 4804 26188 4856 26240
rect 6736 26333 6745 26367
rect 6745 26333 6779 26367
rect 6779 26333 6788 26367
rect 6736 26324 6788 26333
rect 6644 26256 6696 26308
rect 8852 26324 8904 26376
rect 8208 26299 8260 26308
rect 8208 26265 8217 26299
rect 8217 26265 8251 26299
rect 8251 26265 8260 26299
rect 8208 26256 8260 26265
rect 8392 26299 8444 26308
rect 8392 26265 8417 26299
rect 8417 26265 8444 26299
rect 9772 26324 9824 26376
rect 8392 26256 8444 26265
rect 11704 26392 11756 26444
rect 9956 26188 10008 26240
rect 11244 26324 11296 26376
rect 11428 26324 11480 26376
rect 12164 26324 12216 26376
rect 12256 26324 12308 26376
rect 13820 26392 13872 26444
rect 17960 26392 18012 26444
rect 21640 26435 21692 26444
rect 10784 26256 10836 26308
rect 12716 26299 12768 26308
rect 12716 26265 12725 26299
rect 12725 26265 12759 26299
rect 12759 26265 12768 26299
rect 12716 26256 12768 26265
rect 12992 26324 13044 26376
rect 13544 26324 13596 26376
rect 15292 26324 15344 26376
rect 19432 26324 19484 26376
rect 21640 26401 21649 26435
rect 21649 26401 21683 26435
rect 21683 26401 21692 26435
rect 21640 26392 21692 26401
rect 20628 26324 20680 26376
rect 13176 26256 13228 26308
rect 13636 26256 13688 26308
rect 14188 26256 14240 26308
rect 12532 26188 12584 26240
rect 13360 26188 13412 26240
rect 14280 26188 14332 26240
rect 14924 26256 14976 26308
rect 18144 26299 18196 26308
rect 18144 26265 18153 26299
rect 18153 26265 18187 26299
rect 18187 26265 18196 26299
rect 18144 26256 18196 26265
rect 20812 26299 20864 26308
rect 20812 26265 20821 26299
rect 20821 26265 20855 26299
rect 20855 26265 20864 26299
rect 20812 26256 20864 26265
rect 20904 26256 20956 26308
rect 21272 26256 21324 26308
rect 21640 26256 21692 26308
rect 21916 26256 21968 26308
rect 15752 26231 15804 26240
rect 15752 26197 15761 26231
rect 15761 26197 15795 26231
rect 15795 26197 15804 26231
rect 15752 26188 15804 26197
rect 19524 26188 19576 26240
rect 6378 26086 6430 26138
rect 6442 26086 6494 26138
rect 6506 26086 6558 26138
rect 6570 26086 6622 26138
rect 6634 26086 6686 26138
rect 11806 26086 11858 26138
rect 11870 26086 11922 26138
rect 11934 26086 11986 26138
rect 11998 26086 12050 26138
rect 12062 26086 12114 26138
rect 17234 26086 17286 26138
rect 17298 26086 17350 26138
rect 17362 26086 17414 26138
rect 17426 26086 17478 26138
rect 17490 26086 17542 26138
rect 22662 26086 22714 26138
rect 22726 26086 22778 26138
rect 22790 26086 22842 26138
rect 22854 26086 22906 26138
rect 22918 26086 22970 26138
rect 1584 25984 1636 26036
rect 2228 25916 2280 25968
rect 3240 25984 3292 26036
rect 5540 25984 5592 26036
rect 2780 25916 2832 25968
rect 9128 25959 9180 25968
rect 1676 25848 1728 25900
rect 2412 25848 2464 25900
rect 3056 25848 3108 25900
rect 4252 25848 4304 25900
rect 4436 25848 4488 25900
rect 6184 25848 6236 25900
rect 7012 25848 7064 25900
rect 9128 25925 9155 25959
rect 9155 25925 9180 25959
rect 9128 25916 9180 25925
rect 10140 25984 10192 26036
rect 11060 25984 11112 26036
rect 11704 25984 11756 26036
rect 4068 25780 4120 25832
rect 9680 25780 9732 25832
rect 11428 25916 11480 25968
rect 12256 25984 12308 26036
rect 13912 25984 13964 26036
rect 18144 25984 18196 26036
rect 22468 25984 22520 26036
rect 10324 25848 10376 25900
rect 10508 25848 10560 25900
rect 12164 25916 12216 25968
rect 15752 25916 15804 25968
rect 2044 25712 2096 25764
rect 2136 25755 2188 25764
rect 2136 25721 2145 25755
rect 2145 25721 2179 25755
rect 2179 25721 2188 25755
rect 2136 25712 2188 25721
rect 3424 25712 3476 25764
rect 8852 25712 8904 25764
rect 1952 25687 2004 25696
rect 1952 25653 1961 25687
rect 1961 25653 1995 25687
rect 1995 25653 2004 25687
rect 1952 25644 2004 25653
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 3240 25644 3292 25696
rect 3608 25644 3660 25696
rect 7656 25687 7708 25696
rect 7656 25653 7665 25687
rect 7665 25653 7699 25687
rect 7699 25653 7708 25687
rect 7656 25644 7708 25653
rect 9772 25712 9824 25764
rect 13268 25848 13320 25900
rect 14372 25848 14424 25900
rect 19432 25848 19484 25900
rect 19708 25848 19760 25900
rect 20352 25848 20404 25900
rect 13912 25780 13964 25832
rect 19892 25780 19944 25832
rect 21732 25848 21784 25900
rect 21088 25823 21140 25832
rect 21088 25789 21097 25823
rect 21097 25789 21131 25823
rect 21131 25789 21140 25823
rect 21088 25780 21140 25789
rect 14280 25712 14332 25764
rect 22100 25712 22152 25764
rect 11060 25644 11112 25696
rect 11796 25687 11848 25696
rect 11796 25653 11805 25687
rect 11805 25653 11839 25687
rect 11839 25653 11848 25687
rect 11796 25644 11848 25653
rect 12256 25687 12308 25696
rect 12256 25653 12265 25687
rect 12265 25653 12299 25687
rect 12299 25653 12308 25687
rect 12256 25644 12308 25653
rect 12440 25644 12492 25696
rect 13084 25644 13136 25696
rect 13544 25644 13596 25696
rect 20536 25644 20588 25696
rect 21180 25644 21232 25696
rect 21272 25644 21324 25696
rect 22008 25644 22060 25696
rect 3664 25542 3716 25594
rect 3728 25542 3780 25594
rect 3792 25542 3844 25594
rect 3856 25542 3908 25594
rect 3920 25542 3972 25594
rect 9092 25542 9144 25594
rect 9156 25542 9208 25594
rect 9220 25542 9272 25594
rect 9284 25542 9336 25594
rect 9348 25542 9400 25594
rect 14520 25542 14572 25594
rect 14584 25542 14636 25594
rect 14648 25542 14700 25594
rect 14712 25542 14764 25594
rect 14776 25542 14828 25594
rect 19948 25542 20000 25594
rect 20012 25542 20064 25594
rect 20076 25542 20128 25594
rect 20140 25542 20192 25594
rect 20204 25542 20256 25594
rect 1584 25483 1636 25492
rect 1584 25449 1593 25483
rect 1593 25449 1627 25483
rect 1627 25449 1636 25483
rect 1584 25440 1636 25449
rect 2320 25440 2372 25492
rect 6276 25440 6328 25492
rect 7840 25483 7892 25492
rect 7840 25449 7849 25483
rect 7849 25449 7883 25483
rect 7883 25449 7892 25483
rect 7840 25440 7892 25449
rect 11796 25440 11848 25492
rect 13268 25483 13320 25492
rect 4252 25415 4304 25424
rect 4252 25381 4261 25415
rect 4261 25381 4295 25415
rect 4295 25381 4304 25415
rect 4252 25372 4304 25381
rect 4528 25372 4580 25424
rect 7656 25372 7708 25424
rect 13268 25449 13277 25483
rect 13277 25449 13311 25483
rect 13311 25449 13320 25483
rect 13268 25440 13320 25449
rect 19340 25440 19392 25492
rect 19800 25440 19852 25492
rect 9772 25304 9824 25356
rect 12716 25372 12768 25424
rect 20444 25440 20496 25492
rect 20904 25483 20956 25492
rect 20904 25449 20913 25483
rect 20913 25449 20947 25483
rect 20947 25449 20956 25483
rect 20904 25440 20956 25449
rect 20720 25372 20772 25424
rect 2688 25279 2740 25288
rect 2688 25245 2706 25279
rect 2706 25245 2740 25279
rect 2688 25236 2740 25245
rect 4252 25236 4304 25288
rect 5080 25279 5132 25288
rect 5080 25245 5089 25279
rect 5089 25245 5123 25279
rect 5123 25245 5132 25279
rect 5080 25236 5132 25245
rect 6920 25236 6972 25288
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 8484 25236 8536 25288
rect 10324 25236 10376 25288
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 12624 25236 12676 25288
rect 13360 25279 13412 25288
rect 13360 25245 13369 25279
rect 13369 25245 13403 25279
rect 13403 25245 13412 25279
rect 13360 25236 13412 25245
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 20536 25236 20588 25288
rect 22376 25236 22428 25288
rect 2780 25168 2832 25220
rect 4068 25168 4120 25220
rect 2136 25100 2188 25152
rect 5632 25168 5684 25220
rect 11060 25168 11112 25220
rect 13452 25168 13504 25220
rect 21640 25168 21692 25220
rect 4620 25100 4672 25152
rect 4896 25143 4948 25152
rect 4896 25109 4905 25143
rect 4905 25109 4939 25143
rect 4939 25109 4948 25143
rect 4896 25100 4948 25109
rect 10600 25100 10652 25152
rect 10692 25100 10744 25152
rect 11520 25100 11572 25152
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 20076 25100 20128 25152
rect 20536 25100 20588 25152
rect 20628 25100 20680 25152
rect 6378 24998 6430 25050
rect 6442 24998 6494 25050
rect 6506 24998 6558 25050
rect 6570 24998 6622 25050
rect 6634 24998 6686 25050
rect 11806 24998 11858 25050
rect 11870 24998 11922 25050
rect 11934 24998 11986 25050
rect 11998 24998 12050 25050
rect 12062 24998 12114 25050
rect 17234 24998 17286 25050
rect 17298 24998 17350 25050
rect 17362 24998 17414 25050
rect 17426 24998 17478 25050
rect 17490 24998 17542 25050
rect 22662 24998 22714 25050
rect 22726 24998 22778 25050
rect 22790 24998 22842 25050
rect 22854 24998 22906 25050
rect 22918 24998 22970 25050
rect 2044 24896 2096 24948
rect 6184 24896 6236 24948
rect 8852 24896 8904 24948
rect 2320 24828 2372 24880
rect 2780 24828 2832 24880
rect 2688 24803 2740 24812
rect 3424 24828 3476 24880
rect 4804 24828 4856 24880
rect 7104 24828 7156 24880
rect 10508 24828 10560 24880
rect 2688 24769 2706 24803
rect 2706 24769 2740 24803
rect 2688 24760 2740 24769
rect 3608 24803 3660 24812
rect 3608 24769 3627 24803
rect 3627 24769 3660 24803
rect 3608 24760 3660 24769
rect 3332 24692 3384 24744
rect 4068 24760 4120 24812
rect 5080 24760 5132 24812
rect 4988 24692 5040 24744
rect 6276 24760 6328 24812
rect 7472 24760 7524 24812
rect 7564 24760 7616 24812
rect 8300 24760 8352 24812
rect 10968 24896 11020 24948
rect 5264 24624 5316 24676
rect 5356 24667 5408 24676
rect 5356 24633 5365 24667
rect 5365 24633 5399 24667
rect 5399 24633 5408 24667
rect 5356 24624 5408 24633
rect 9680 24624 9732 24676
rect 9864 24624 9916 24676
rect 10692 24692 10744 24744
rect 11612 24760 11664 24812
rect 14280 24828 14332 24880
rect 19340 24828 19392 24880
rect 12808 24803 12860 24812
rect 12808 24769 12817 24803
rect 12817 24769 12851 24803
rect 12851 24769 12860 24803
rect 12808 24760 12860 24769
rect 17408 24760 17460 24812
rect 17040 24692 17092 24744
rect 18052 24692 18104 24744
rect 21088 24896 21140 24948
rect 21640 24896 21692 24948
rect 20168 24828 20220 24880
rect 20996 24828 21048 24880
rect 21548 24760 21600 24812
rect 22100 24760 22152 24812
rect 22376 24692 22428 24744
rect 19800 24624 19852 24676
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2780 24556 2832 24608
rect 3608 24556 3660 24608
rect 4160 24556 4212 24608
rect 4252 24556 4304 24608
rect 4344 24556 4396 24608
rect 4528 24556 4580 24608
rect 5080 24556 5132 24608
rect 8576 24599 8628 24608
rect 8576 24565 8585 24599
rect 8585 24565 8619 24599
rect 8619 24565 8628 24599
rect 8576 24556 8628 24565
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 10508 24556 10560 24608
rect 10692 24556 10744 24608
rect 17776 24556 17828 24608
rect 18696 24599 18748 24608
rect 18696 24565 18705 24599
rect 18705 24565 18739 24599
rect 18739 24565 18748 24599
rect 18696 24556 18748 24565
rect 19616 24599 19668 24608
rect 19616 24565 19625 24599
rect 19625 24565 19659 24599
rect 19659 24565 19668 24599
rect 19616 24556 19668 24565
rect 21456 24556 21508 24608
rect 3664 24454 3716 24506
rect 3728 24454 3780 24506
rect 3792 24454 3844 24506
rect 3856 24454 3908 24506
rect 3920 24454 3972 24506
rect 9092 24454 9144 24506
rect 9156 24454 9208 24506
rect 9220 24454 9272 24506
rect 9284 24454 9336 24506
rect 9348 24454 9400 24506
rect 14520 24454 14572 24506
rect 14584 24454 14636 24506
rect 14648 24454 14700 24506
rect 14712 24454 14764 24506
rect 14776 24454 14828 24506
rect 19948 24454 20000 24506
rect 20012 24454 20064 24506
rect 20076 24454 20128 24506
rect 20140 24454 20192 24506
rect 20204 24454 20256 24506
rect 1676 24352 1728 24404
rect 4252 24352 4304 24404
rect 4436 24352 4488 24404
rect 5448 24352 5500 24404
rect 9588 24395 9640 24404
rect 9588 24361 9597 24395
rect 9597 24361 9631 24395
rect 9631 24361 9640 24395
rect 9588 24352 9640 24361
rect 10416 24395 10468 24404
rect 10416 24361 10425 24395
rect 10425 24361 10459 24395
rect 10459 24361 10468 24395
rect 10416 24352 10468 24361
rect 11152 24352 11204 24404
rect 17408 24395 17460 24404
rect 17408 24361 17417 24395
rect 17417 24361 17451 24395
rect 17451 24361 17460 24395
rect 17408 24352 17460 24361
rect 17592 24352 17644 24404
rect 19432 24352 19484 24404
rect 19616 24352 19668 24404
rect 20720 24352 20772 24404
rect 21916 24352 21968 24404
rect 6644 24327 6696 24336
rect 4712 24216 4764 24268
rect 5448 24216 5500 24268
rect 2688 24191 2740 24200
rect 2688 24157 2706 24191
rect 2706 24157 2740 24191
rect 2688 24148 2740 24157
rect 2320 24080 2372 24132
rect 3608 24148 3660 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 3424 24080 3476 24132
rect 5080 24148 5132 24200
rect 4436 24080 4488 24132
rect 5356 24123 5408 24132
rect 5356 24089 5365 24123
rect 5365 24089 5399 24123
rect 5399 24089 5408 24123
rect 5356 24080 5408 24089
rect 6644 24293 6653 24327
rect 6653 24293 6687 24327
rect 6687 24293 6696 24327
rect 6644 24284 6696 24293
rect 7196 24284 7248 24336
rect 7472 24284 7524 24336
rect 8576 24284 8628 24336
rect 13176 24284 13228 24336
rect 21272 24284 21324 24336
rect 10048 24216 10100 24268
rect 12348 24216 12400 24268
rect 5632 24148 5684 24200
rect 9496 24148 9548 24200
rect 11336 24148 11388 24200
rect 19340 24216 19392 24268
rect 17684 24148 17736 24200
rect 6184 24123 6236 24132
rect 6184 24089 6193 24123
rect 6193 24089 6227 24123
rect 6227 24089 6236 24123
rect 6184 24080 6236 24089
rect 11428 24080 11480 24132
rect 19064 24148 19116 24200
rect 19248 24148 19300 24200
rect 19616 24148 19668 24200
rect 19984 24148 20036 24200
rect 22008 24191 22060 24200
rect 22008 24157 22026 24191
rect 22026 24157 22060 24191
rect 22008 24148 22060 24157
rect 22376 24148 22428 24200
rect 1676 24012 1728 24064
rect 2504 24012 2556 24064
rect 5172 24055 5224 24064
rect 5172 24021 5199 24055
rect 5199 24021 5224 24055
rect 5172 24012 5224 24021
rect 5816 24055 5868 24064
rect 5816 24021 5825 24055
rect 5825 24021 5859 24055
rect 5859 24021 5868 24055
rect 5816 24012 5868 24021
rect 17868 24012 17920 24064
rect 19984 24012 20036 24064
rect 22192 24080 22244 24132
rect 6378 23910 6430 23962
rect 6442 23910 6494 23962
rect 6506 23910 6558 23962
rect 6570 23910 6622 23962
rect 6634 23910 6686 23962
rect 11806 23910 11858 23962
rect 11870 23910 11922 23962
rect 11934 23910 11986 23962
rect 11998 23910 12050 23962
rect 12062 23910 12114 23962
rect 17234 23910 17286 23962
rect 17298 23910 17350 23962
rect 17362 23910 17414 23962
rect 17426 23910 17478 23962
rect 17490 23910 17542 23962
rect 22662 23910 22714 23962
rect 22726 23910 22778 23962
rect 22790 23910 22842 23962
rect 22854 23910 22906 23962
rect 22918 23910 22970 23962
rect 3148 23808 3200 23860
rect 4068 23808 4120 23860
rect 4160 23808 4212 23860
rect 6184 23808 6236 23860
rect 10876 23808 10928 23860
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 1584 23715 1636 23724
rect 1584 23681 1593 23715
rect 1593 23681 1627 23715
rect 1627 23681 1636 23715
rect 1584 23672 1636 23681
rect 2228 23672 2280 23724
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 4712 23740 4764 23792
rect 5080 23740 5132 23792
rect 5356 23740 5408 23792
rect 8116 23783 8168 23792
rect 2596 23647 2648 23656
rect 2596 23613 2605 23647
rect 2605 23613 2639 23647
rect 2639 23613 2648 23647
rect 2596 23604 2648 23613
rect 3148 23468 3200 23520
rect 4436 23672 4488 23724
rect 5908 23715 5960 23724
rect 5908 23681 5917 23715
rect 5917 23681 5951 23715
rect 5951 23681 5960 23715
rect 6736 23715 6788 23724
rect 5908 23672 5960 23681
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 8116 23749 8125 23783
rect 8125 23749 8159 23783
rect 8159 23749 8168 23783
rect 8116 23740 8168 23749
rect 12348 23740 12400 23792
rect 16672 23740 16724 23792
rect 17868 23740 17920 23792
rect 19340 23808 19392 23860
rect 20444 23808 20496 23860
rect 20720 23808 20772 23860
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 5356 23604 5408 23656
rect 5448 23536 5500 23588
rect 11244 23672 11296 23724
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 19064 23715 19116 23724
rect 19064 23681 19073 23715
rect 19073 23681 19107 23715
rect 19107 23681 19116 23715
rect 19064 23672 19116 23681
rect 19340 23715 19392 23724
rect 19340 23681 19349 23715
rect 19349 23681 19383 23715
rect 19383 23681 19392 23715
rect 19340 23672 19392 23681
rect 19524 23672 19576 23724
rect 21364 23672 21416 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 21548 23604 21600 23656
rect 22376 23604 22428 23656
rect 19432 23536 19484 23588
rect 5356 23468 5408 23520
rect 6828 23468 6880 23520
rect 18604 23511 18656 23520
rect 18604 23477 18613 23511
rect 18613 23477 18647 23511
rect 18647 23477 18656 23511
rect 18604 23468 18656 23477
rect 20444 23468 20496 23520
rect 21272 23468 21324 23520
rect 3664 23366 3716 23418
rect 3728 23366 3780 23418
rect 3792 23366 3844 23418
rect 3856 23366 3908 23418
rect 3920 23366 3972 23418
rect 9092 23366 9144 23418
rect 9156 23366 9208 23418
rect 9220 23366 9272 23418
rect 9284 23366 9336 23418
rect 9348 23366 9400 23418
rect 14520 23366 14572 23418
rect 14584 23366 14636 23418
rect 14648 23366 14700 23418
rect 14712 23366 14764 23418
rect 14776 23366 14828 23418
rect 19948 23366 20000 23418
rect 20012 23366 20064 23418
rect 20076 23366 20128 23418
rect 20140 23366 20192 23418
rect 20204 23366 20256 23418
rect 3424 23264 3476 23316
rect 5908 23307 5960 23316
rect 5908 23273 5917 23307
rect 5917 23273 5951 23307
rect 5951 23273 5960 23307
rect 5908 23264 5960 23273
rect 6092 23264 6144 23316
rect 9864 23264 9916 23316
rect 16856 23307 16908 23316
rect 16856 23273 16865 23307
rect 16865 23273 16899 23307
rect 16899 23273 16908 23307
rect 16856 23264 16908 23273
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 4896 23196 4948 23248
rect 6920 23196 6972 23248
rect 17040 23239 17092 23248
rect 17040 23205 17049 23239
rect 17049 23205 17083 23239
rect 17083 23205 17092 23239
rect 17040 23196 17092 23205
rect 17868 23239 17920 23248
rect 17868 23205 17877 23239
rect 17877 23205 17911 23239
rect 17911 23205 17920 23239
rect 17868 23196 17920 23205
rect 19432 23264 19484 23316
rect 20352 23264 20404 23316
rect 20904 23264 20956 23316
rect 22100 23196 22152 23248
rect 2964 23128 3016 23180
rect 2872 23060 2924 23112
rect 3148 23060 3200 23112
rect 4160 23103 4212 23112
rect 4160 23069 4164 23103
rect 4164 23069 4198 23103
rect 4198 23069 4212 23103
rect 4160 23060 4212 23069
rect 2964 22992 3016 23044
rect 4068 22992 4120 23044
rect 4620 23103 4672 23112
rect 4620 23069 4629 23103
rect 4629 23069 4663 23103
rect 4663 23069 4672 23103
rect 5356 23128 5408 23180
rect 18236 23128 18288 23180
rect 20076 23128 20128 23180
rect 20628 23128 20680 23180
rect 21088 23128 21140 23180
rect 21364 23128 21416 23180
rect 4620 23060 4672 23069
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 19616 23060 19668 23112
rect 19892 23060 19944 23112
rect 20444 23103 20496 23112
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 22284 23060 22336 23112
rect 4804 22992 4856 23044
rect 5448 23035 5500 23044
rect 5448 23001 5457 23035
rect 5457 23001 5491 23035
rect 5491 23001 5500 23035
rect 5448 22992 5500 23001
rect 16672 23035 16724 23044
rect 16672 23001 16681 23035
rect 16681 23001 16715 23035
rect 16715 23001 16724 23035
rect 16672 22992 16724 23001
rect 17224 22992 17276 23044
rect 3148 22924 3200 22976
rect 4620 22924 4672 22976
rect 5172 22924 5224 22976
rect 18328 22992 18380 23044
rect 19064 22992 19116 23044
rect 20904 22992 20956 23044
rect 17684 22924 17736 22976
rect 19524 22924 19576 22976
rect 19800 22967 19852 22976
rect 19800 22933 19809 22967
rect 19809 22933 19843 22967
rect 19843 22933 19852 22967
rect 19800 22924 19852 22933
rect 21272 22924 21324 22976
rect 6378 22822 6430 22874
rect 6442 22822 6494 22874
rect 6506 22822 6558 22874
rect 6570 22822 6622 22874
rect 6634 22822 6686 22874
rect 11806 22822 11858 22874
rect 11870 22822 11922 22874
rect 11934 22822 11986 22874
rect 11998 22822 12050 22874
rect 12062 22822 12114 22874
rect 17234 22822 17286 22874
rect 17298 22822 17350 22874
rect 17362 22822 17414 22874
rect 17426 22822 17478 22874
rect 17490 22822 17542 22874
rect 22662 22822 22714 22874
rect 22726 22822 22778 22874
rect 22790 22822 22842 22874
rect 22854 22822 22906 22874
rect 22918 22822 22970 22874
rect 5172 22720 5224 22772
rect 7104 22763 7156 22772
rect 7104 22729 7113 22763
rect 7113 22729 7147 22763
rect 7147 22729 7156 22763
rect 7104 22720 7156 22729
rect 18236 22763 18288 22772
rect 18236 22729 18245 22763
rect 18245 22729 18279 22763
rect 18279 22729 18288 22763
rect 18236 22720 18288 22729
rect 19294 22720 19346 22772
rect 19708 22720 19760 22772
rect 20076 22763 20128 22772
rect 3424 22652 3476 22704
rect 6828 22652 6880 22704
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2320 22584 2372 22636
rect 4068 22584 4120 22636
rect 6092 22584 6144 22636
rect 2688 22516 2740 22568
rect 5356 22516 5408 22568
rect 8116 22584 8168 22636
rect 17868 22516 17920 22568
rect 18696 22584 18748 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19432 22652 19484 22704
rect 20076 22729 20085 22763
rect 20085 22729 20119 22763
rect 20119 22729 20128 22763
rect 20076 22720 20128 22729
rect 20168 22720 20220 22772
rect 21640 22720 21692 22772
rect 20720 22652 20772 22704
rect 21456 22652 21508 22704
rect 20168 22584 20220 22636
rect 2320 22380 2372 22432
rect 2872 22448 2924 22500
rect 3884 22448 3936 22500
rect 3056 22380 3108 22432
rect 4160 22380 4212 22432
rect 4620 22423 4672 22432
rect 4620 22389 4629 22423
rect 4629 22389 4663 22423
rect 4663 22389 4672 22423
rect 4620 22380 4672 22389
rect 6736 22448 6788 22500
rect 21824 22584 21876 22636
rect 21548 22516 21600 22568
rect 22100 22584 22152 22636
rect 17592 22423 17644 22432
rect 17592 22389 17601 22423
rect 17601 22389 17635 22423
rect 17635 22389 17644 22423
rect 17592 22380 17644 22389
rect 18880 22380 18932 22432
rect 19616 22380 19668 22432
rect 20076 22380 20128 22432
rect 21916 22380 21968 22432
rect 3664 22278 3716 22330
rect 3728 22278 3780 22330
rect 3792 22278 3844 22330
rect 3856 22278 3908 22330
rect 3920 22278 3972 22330
rect 9092 22278 9144 22330
rect 9156 22278 9208 22330
rect 9220 22278 9272 22330
rect 9284 22278 9336 22330
rect 9348 22278 9400 22330
rect 14520 22278 14572 22330
rect 14584 22278 14636 22330
rect 14648 22278 14700 22330
rect 14712 22278 14764 22330
rect 14776 22278 14828 22330
rect 19948 22278 20000 22330
rect 20012 22278 20064 22330
rect 20076 22278 20128 22330
rect 20140 22278 20192 22330
rect 20204 22278 20256 22330
rect 2228 22176 2280 22228
rect 3424 22176 3476 22228
rect 4620 22176 4672 22228
rect 5356 22176 5408 22228
rect 20812 22176 20864 22228
rect 4988 22108 5040 22160
rect 16856 22108 16908 22160
rect 19340 22108 19392 22160
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 4068 22040 4120 22092
rect 4252 22040 4304 22092
rect 4712 22040 4764 22092
rect 7288 22040 7340 22092
rect 10600 22083 10652 22092
rect 10600 22049 10609 22083
rect 10609 22049 10643 22083
rect 10643 22049 10652 22083
rect 10600 22040 10652 22049
rect 21088 22108 21140 22160
rect 1860 22015 1912 22024
rect 1860 21981 1894 22015
rect 1894 21981 1912 22015
rect 1860 21972 1912 21981
rect 2412 21972 2464 22024
rect 3884 21972 3936 22024
rect 4804 22015 4856 22024
rect 2872 21904 2924 21956
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 5632 21972 5684 22024
rect 11704 21972 11756 22024
rect 18604 22015 18656 22024
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 17684 21904 17736 21956
rect 19340 21972 19392 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 21272 22040 21324 22092
rect 19984 21904 20036 21956
rect 21180 21972 21232 22024
rect 2504 21836 2556 21888
rect 10416 21836 10468 21888
rect 17776 21836 17828 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 18788 21836 18840 21845
rect 20260 21879 20312 21888
rect 20260 21845 20269 21879
rect 20269 21845 20303 21879
rect 20303 21845 20312 21879
rect 20260 21836 20312 21845
rect 20720 21904 20772 21956
rect 21548 21904 21600 21956
rect 20536 21836 20588 21888
rect 21088 21836 21140 21888
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 2136 21675 2188 21684
rect 2136 21641 2145 21675
rect 2145 21641 2179 21675
rect 2179 21641 2188 21675
rect 2136 21632 2188 21641
rect 2596 21675 2648 21684
rect 2596 21641 2605 21675
rect 2605 21641 2639 21675
rect 2639 21641 2648 21675
rect 2596 21632 2648 21641
rect 3148 21632 3200 21684
rect 4436 21632 4488 21684
rect 4896 21675 4948 21684
rect 4896 21641 4905 21675
rect 4905 21641 4939 21675
rect 4939 21641 4948 21675
rect 5356 21675 5408 21684
rect 4896 21632 4948 21641
rect 5356 21641 5365 21675
rect 5365 21641 5399 21675
rect 5399 21641 5408 21675
rect 5356 21632 5408 21641
rect 18788 21632 18840 21684
rect 2228 21564 2280 21616
rect 19432 21564 19484 21616
rect 20260 21564 20312 21616
rect 20536 21564 20588 21616
rect 20720 21564 20772 21616
rect 21272 21632 21324 21684
rect 21088 21607 21140 21616
rect 21088 21573 21097 21607
rect 21097 21573 21131 21607
rect 21131 21573 21140 21607
rect 21088 21564 21140 21573
rect 22192 21564 22244 21616
rect 2412 21496 2464 21548
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 4160 21539 4212 21548
rect 2136 21428 2188 21480
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 9864 21496 9916 21548
rect 10600 21539 10652 21548
rect 10600 21505 10609 21539
rect 10609 21505 10643 21539
rect 10643 21505 10652 21539
rect 10600 21496 10652 21505
rect 20812 21496 20864 21548
rect 3148 21428 3200 21480
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 19524 21428 19576 21480
rect 19984 21428 20036 21480
rect 20720 21428 20772 21480
rect 5816 21360 5868 21412
rect 19616 21360 19668 21412
rect 10324 21292 10376 21344
rect 17776 21292 17828 21344
rect 19248 21292 19300 21344
rect 21272 21539 21324 21548
rect 21272 21505 21317 21539
rect 21317 21505 21324 21539
rect 21272 21496 21324 21505
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22008 21292 22060 21344
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 2136 21131 2188 21140
rect 2136 21097 2145 21131
rect 2145 21097 2179 21131
rect 2179 21097 2188 21131
rect 2136 21088 2188 21097
rect 3240 21088 3292 21140
rect 4896 21088 4948 21140
rect 11704 21131 11756 21140
rect 11704 21097 11713 21131
rect 11713 21097 11747 21131
rect 11747 21097 11756 21131
rect 11704 21088 11756 21097
rect 19524 21088 19576 21140
rect 20628 21088 20680 21140
rect 1768 21020 1820 21072
rect 3332 20952 3384 21004
rect 4620 20952 4672 21004
rect 7380 20952 7432 21004
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 17776 20952 17828 21004
rect 21548 21088 21600 21140
rect 22284 21131 22336 21140
rect 22284 21097 22293 21131
rect 22293 21097 22327 21131
rect 22327 21097 22336 21131
rect 22284 21088 22336 21097
rect 1768 20884 1820 20936
rect 4160 20884 4212 20936
rect 2872 20816 2924 20868
rect 8760 20884 8812 20936
rect 10416 20884 10468 20936
rect 19708 20884 19760 20936
rect 20996 20884 21048 20936
rect 19800 20816 19852 20868
rect 21640 20816 21692 20868
rect 3424 20748 3476 20800
rect 7104 20791 7156 20800
rect 7104 20757 7113 20791
rect 7113 20757 7147 20791
rect 7147 20757 7156 20791
rect 7104 20748 7156 20757
rect 18328 20748 18380 20800
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 1952 20544 2004 20596
rect 4804 20544 4856 20596
rect 1768 20519 1820 20528
rect 1768 20485 1777 20519
rect 1777 20485 1811 20519
rect 1811 20485 1820 20519
rect 1768 20476 1820 20485
rect 7104 20476 7156 20528
rect 20904 20544 20956 20596
rect 21732 20544 21784 20596
rect 20536 20476 20588 20528
rect 2320 20408 2372 20460
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 7380 20451 7432 20460
rect 7380 20417 7389 20451
rect 7389 20417 7423 20451
rect 7423 20417 7432 20451
rect 7380 20408 7432 20417
rect 10600 20272 10652 20324
rect 13360 20408 13412 20460
rect 20352 20408 20404 20460
rect 20444 20408 20496 20460
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 8760 20247 8812 20256
rect 8760 20213 8769 20247
rect 8769 20213 8803 20247
rect 8803 20213 8812 20247
rect 8760 20204 8812 20213
rect 12532 20204 12584 20256
rect 16856 20340 16908 20392
rect 14280 20204 14332 20256
rect 17776 20204 17828 20256
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 22284 20247 22336 20256
rect 22284 20213 22293 20247
rect 22293 20213 22327 20247
rect 22327 20213 22336 20247
rect 22284 20204 22336 20213
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 20812 20000 20864 20052
rect 21916 20043 21968 20052
rect 21916 20009 21925 20043
rect 21925 20009 21959 20043
rect 21959 20009 21968 20043
rect 21916 20000 21968 20009
rect 22192 20000 22244 20052
rect 19616 19864 19668 19916
rect 1492 19796 1544 19848
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 3424 19660 3476 19712
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 1860 19456 1912 19508
rect 11704 19456 11756 19508
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 12394 19320 12446 19372
rect 12532 19363 12584 19372
rect 12532 19329 12550 19363
rect 12550 19329 12584 19363
rect 12532 19320 12584 19329
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 22008 19320 22060 19372
rect 9496 19252 9548 19304
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2780 19116 2832 19168
rect 10968 19159 11020 19168
rect 10968 19125 10977 19159
rect 10977 19125 11011 19159
rect 11011 19125 11020 19159
rect 10968 19116 11020 19125
rect 12256 19116 12308 19168
rect 22192 19116 22244 19168
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 3056 18912 3108 18964
rect 21548 18955 21600 18964
rect 21548 18921 21557 18955
rect 21557 18921 21591 18955
rect 21591 18921 21600 18955
rect 21548 18912 21600 18921
rect 5724 18844 5776 18896
rect 6736 18776 6788 18828
rect 2780 18708 2832 18760
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 9496 18708 9548 18760
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 4620 18640 4672 18692
rect 2872 18572 2924 18624
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 3332 18368 3384 18420
rect 9496 18368 9548 18420
rect 2228 18300 2280 18352
rect 7380 18300 7432 18352
rect 2964 18275 3016 18284
rect 2320 18164 2372 18216
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 7472 18232 7524 18284
rect 3332 18164 3384 18216
rect 2044 18096 2096 18148
rect 22284 18139 22336 18148
rect 22284 18105 22293 18139
rect 22293 18105 22327 18139
rect 22327 18105 22336 18139
rect 22284 18096 22336 18105
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 22192 17824 22244 17876
rect 1492 17620 1544 17672
rect 2596 17620 2648 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 1676 17552 1728 17604
rect 3240 17552 3292 17604
rect 5816 17552 5868 17604
rect 2688 17484 2740 17536
rect 4344 17527 4396 17536
rect 4344 17493 4353 17527
rect 4353 17493 4387 17527
rect 4387 17493 4396 17527
rect 4344 17484 4396 17493
rect 4436 17484 4488 17536
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 5172 17280 5224 17332
rect 4436 17212 4488 17264
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 3516 17144 3568 17196
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 3148 17076 3200 17128
rect 2964 17008 3016 17060
rect 4160 17008 4212 17060
rect 22284 17051 22336 17060
rect 22284 17017 22293 17051
rect 22293 17017 22327 17051
rect 22327 17017 22336 17051
rect 22284 17008 22336 17017
rect 4068 16940 4120 16992
rect 4252 16940 4304 16992
rect 4896 16940 4948 16992
rect 7472 16940 7524 16992
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 1584 16736 1636 16788
rect 2964 16736 3016 16788
rect 4344 16779 4396 16788
rect 3424 16600 3476 16652
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 6000 16779 6052 16788
rect 6000 16745 6009 16779
rect 6009 16745 6043 16779
rect 6043 16745 6052 16779
rect 6000 16736 6052 16745
rect 6092 16668 6144 16720
rect 4896 16600 4948 16652
rect 1860 16575 1912 16584
rect 1860 16541 1894 16575
rect 1894 16541 1912 16575
rect 1860 16532 1912 16541
rect 2228 16532 2280 16584
rect 4344 16532 4396 16584
rect 5540 16532 5592 16584
rect 6000 16532 6052 16584
rect 22008 16600 22060 16652
rect 5172 16507 5224 16516
rect 5172 16473 5181 16507
rect 5181 16473 5215 16507
rect 5215 16473 5224 16507
rect 5172 16464 5224 16473
rect 3056 16396 3108 16448
rect 4344 16439 4396 16448
rect 4344 16405 4353 16439
rect 4353 16405 4387 16439
rect 4387 16405 4396 16439
rect 4344 16396 4396 16405
rect 4804 16396 4856 16448
rect 5264 16396 5316 16448
rect 5816 16439 5868 16448
rect 5816 16405 5825 16439
rect 5825 16405 5859 16439
rect 5859 16405 5868 16439
rect 5816 16396 5868 16405
rect 6000 16439 6052 16448
rect 6000 16405 6027 16439
rect 6027 16405 6052 16439
rect 6000 16396 6052 16405
rect 6276 16396 6328 16448
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 2596 16192 2648 16244
rect 3332 16192 3384 16244
rect 6000 16192 6052 16244
rect 22100 16192 22152 16244
rect 5908 16124 5960 16176
rect 6184 16124 6236 16176
rect 6920 16167 6972 16176
rect 6920 16133 6929 16167
rect 6929 16133 6963 16167
rect 6963 16133 6972 16167
rect 6920 16124 6972 16133
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 2964 16056 3016 16065
rect 6552 16056 6604 16108
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 4896 15988 4948 16040
rect 5540 15988 5592 16040
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 4160 15852 4212 15904
rect 5540 15852 5592 15904
rect 6736 15895 6788 15904
rect 6736 15861 6745 15895
rect 6745 15861 6779 15895
rect 6779 15861 6788 15895
rect 6736 15852 6788 15861
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 2780 15648 2832 15700
rect 3240 15648 3292 15700
rect 4712 15648 4764 15700
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 5908 15691 5960 15700
rect 5908 15657 5917 15691
rect 5917 15657 5951 15691
rect 5951 15657 5960 15691
rect 5908 15648 5960 15657
rect 6552 15691 6604 15700
rect 6552 15657 6561 15691
rect 6561 15657 6595 15691
rect 6595 15657 6604 15691
rect 6552 15648 6604 15657
rect 4252 15580 4304 15632
rect 4804 15580 4856 15632
rect 2964 15512 3016 15564
rect 3240 15512 3292 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 3056 15487 3108 15496
rect 1768 15376 1820 15428
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 4160 15512 4212 15564
rect 4068 15487 4120 15496
rect 4068 15453 4078 15487
rect 4078 15453 4112 15487
rect 4112 15453 4120 15487
rect 4620 15512 4672 15564
rect 4068 15444 4120 15453
rect 4528 15444 4580 15496
rect 2964 15376 3016 15428
rect 3332 15376 3384 15428
rect 6276 15512 6328 15564
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6736 15580 6788 15632
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 10968 15444 11020 15496
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 1952 15308 2004 15360
rect 2228 15308 2280 15360
rect 2320 15308 2372 15360
rect 3608 15308 3660 15360
rect 6184 15308 6236 15360
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 3516 15104 3568 15156
rect 4988 15104 5040 15156
rect 2596 15036 2648 15088
rect 3332 14900 3384 14952
rect 3516 14900 3568 14952
rect 2596 14764 2648 14816
rect 4068 14968 4120 15020
rect 5172 14968 5224 15020
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 4160 14900 4212 14952
rect 4804 14875 4856 14884
rect 4804 14841 4813 14875
rect 4813 14841 4847 14875
rect 4847 14841 4856 14875
rect 4804 14832 4856 14841
rect 22284 14875 22336 14884
rect 22284 14841 22293 14875
rect 22293 14841 22327 14875
rect 22327 14841 22336 14875
rect 22284 14832 22336 14841
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 3976 14560 4028 14612
rect 3240 14492 3292 14544
rect 3700 14424 3752 14476
rect 4344 14467 4396 14476
rect 4344 14433 4353 14467
rect 4353 14433 4387 14467
rect 4387 14433 4396 14467
rect 4344 14424 4396 14433
rect 2872 14356 2924 14408
rect 3884 14356 3936 14408
rect 3424 14288 3476 14340
rect 4160 14331 4212 14340
rect 4160 14297 4169 14331
rect 4169 14297 4203 14331
rect 4203 14297 4212 14331
rect 4160 14288 4212 14297
rect 4804 14288 4856 14340
rect 2688 14220 2740 14272
rect 4620 14220 4672 14272
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 2964 14016 3016 14068
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 2504 13812 2556 13864
rect 3332 13880 3384 13932
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 4252 13880 4304 13932
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 6736 13812 6788 13864
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 2780 13744 2832 13796
rect 3148 13744 3200 13796
rect 2044 13676 2096 13728
rect 2872 13676 2924 13728
rect 3792 13676 3844 13728
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 1768 13472 1820 13524
rect 2412 13472 2464 13524
rect 2688 13472 2740 13524
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 2872 13336 2924 13388
rect 1952 13268 2004 13277
rect 2320 13200 2372 13252
rect 3332 13472 3384 13524
rect 4436 13472 4488 13524
rect 3516 13268 3568 13320
rect 22284 13311 22336 13320
rect 22284 13277 22293 13311
rect 22293 13277 22327 13311
rect 22327 13277 22336 13311
rect 22284 13268 22336 13277
rect 2412 13132 2464 13184
rect 3148 13132 3200 13184
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 4620 12928 4672 12980
rect 3148 12860 3200 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 2872 12792 2924 12844
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3516 12792 3568 12844
rect 3424 12724 3476 12776
rect 2320 12656 2372 12708
rect 2596 12656 2648 12708
rect 3148 12588 3200 12640
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 1676 12384 1728 12436
rect 2780 12384 2832 12436
rect 1952 12316 2004 12368
rect 4068 12384 4120 12436
rect 3240 12248 3292 12300
rect 2780 12180 2832 12232
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 2504 11840 2556 11892
rect 3148 11772 3200 11824
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 22284 11611 22336 11620
rect 22284 11577 22293 11611
rect 22293 11577 22327 11611
rect 22327 11577 22336 11611
rect 22284 11568 22336 11577
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 1768 11296 1820 11348
rect 1492 11092 1544 11144
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 2780 10752 2832 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 22284 10523 22336 10532
rect 22284 10489 22293 10523
rect 22293 10489 22327 10523
rect 22327 10489 22336 10523
rect 22284 10480 22336 10489
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 1492 9120 1544 9172
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 22284 8347 22336 8356
rect 22284 8313 22293 8347
rect 22293 8313 22327 8347
rect 22327 8313 22336 8347
rect 22284 8304 22336 8313
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 22284 7259 22336 7268
rect 22284 7225 22293 7259
rect 22293 7225 22327 7259
rect 22327 7225 22336 7259
rect 22284 7216 22336 7225
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 22284 6783 22336 6792
rect 22284 6749 22293 6783
rect 22293 6749 22327 6783
rect 22327 6749 22336 6783
rect 22284 6740 22336 6749
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 7472 6264 7524 6316
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 22284 5083 22336 5092
rect 22284 5049 22293 5083
rect 22293 5049 22327 5083
rect 22327 5049 22336 5083
rect 22284 5040 22336 5049
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 22284 3995 22336 4004
rect 22284 3961 22293 3995
rect 22293 3961 22327 3995
rect 22327 3961 22336 3995
rect 22284 3952 22336 3961
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 22284 3519 22336 3528
rect 22284 3485 22293 3519
rect 22293 3485 22327 3519
rect 22327 3485 22336 3519
rect 22284 3476 22336 3485
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 1400 2796 1452 2848
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 1214 29200 1270 30000
rect 2042 29322 2098 30000
rect 2870 29322 2926 30000
rect 2042 29294 2360 29322
rect 2042 29200 2098 29294
rect 1228 25401 1256 29200
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1584 27056 1636 27062
rect 1584 26998 1636 27004
rect 1596 26314 1624 26998
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 26042 1624 26250
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1596 25498 1624 25978
rect 1688 25906 1716 26726
rect 1676 25900 1728 25906
rect 1676 25842 1728 25848
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 1214 25392 1270 25401
rect 1214 25327 1270 25336
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1596 23730 1624 24550
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1688 24070 1716 24346
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1584 23724 1636 23730
rect 1584 23666 1636 23672
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1596 22642 1624 23054
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1596 22098 1624 22578
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1688 20890 1716 24006
rect 1780 21078 1808 27406
rect 1860 27328 1912 27334
rect 1860 27270 1912 27276
rect 1872 22030 1900 27270
rect 2044 26988 2096 26994
rect 2044 26930 2096 26936
rect 2056 26586 2084 26930
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 2228 26512 2280 26518
rect 2228 26454 2280 26460
rect 2240 25974 2268 26454
rect 2228 25968 2280 25974
rect 2228 25910 2280 25916
rect 2044 25764 2096 25770
rect 2044 25706 2096 25712
rect 2136 25764 2188 25770
rect 2136 25706 2188 25712
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1768 21072 1820 21078
rect 1768 21014 1820 21020
rect 1768 20936 1820 20942
rect 1688 20884 1768 20890
rect 1688 20878 1820 20884
rect 1688 20862 1808 20878
rect 1780 20534 1808 20862
rect 1964 20602 1992 25638
rect 2056 24954 2084 25706
rect 2148 25158 2176 25706
rect 2136 25152 2188 25158
rect 2136 25094 2188 25100
rect 2044 24948 2096 24954
rect 2044 24890 2096 24896
rect 2240 23730 2268 25910
rect 2332 25498 2360 29294
rect 2870 29294 3188 29322
rect 2870 29200 2926 29294
rect 2412 27328 2464 27334
rect 2412 27270 2464 27276
rect 2964 27328 3016 27334
rect 2964 27270 3016 27276
rect 2424 26382 2452 27270
rect 2504 26784 2556 26790
rect 2688 26784 2740 26790
rect 2556 26744 2636 26772
rect 2504 26726 2556 26732
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 2504 26308 2556 26314
rect 2504 26250 2556 26256
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2320 25492 2372 25498
rect 2320 25434 2372 25440
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2332 24138 2360 24822
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2240 22234 2268 23666
rect 2332 22642 2360 24074
rect 2424 23610 2452 25842
rect 2516 24857 2544 26250
rect 2502 24848 2558 24857
rect 2502 24783 2558 24792
rect 2504 24064 2556 24070
rect 2608 24041 2636 26744
rect 2688 26726 2740 26732
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2700 25294 2728 26726
rect 2780 26512 2832 26518
rect 2780 26454 2832 26460
rect 2792 25974 2820 26454
rect 2780 25968 2832 25974
rect 2780 25910 2832 25916
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2780 25220 2832 25226
rect 2780 25162 2832 25168
rect 2792 24886 2820 25162
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2700 24721 2728 24754
rect 2686 24712 2742 24721
rect 2686 24647 2742 24656
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2686 24304 2742 24313
rect 2686 24239 2742 24248
rect 2700 24206 2728 24239
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2504 24006 2556 24012
rect 2594 24032 2650 24041
rect 2516 23730 2544 24006
rect 2594 23967 2650 23976
rect 2608 23746 2636 23967
rect 2504 23724 2556 23730
rect 2608 23718 2728 23746
rect 2504 23666 2556 23672
rect 2596 23656 2648 23662
rect 2424 23582 2544 23610
rect 2596 23598 2648 23604
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2320 22432 2372 22438
rect 2320 22374 2372 22380
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2134 21720 2190 21729
rect 2134 21655 2136 21664
rect 2188 21655 2190 21664
rect 2136 21626 2188 21632
rect 2240 21622 2268 22170
rect 2228 21616 2280 21622
rect 2228 21558 2280 21564
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2148 21146 2176 21422
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1768 20528 1820 20534
rect 1768 20470 1820 20476
rect 2332 20466 2360 22374
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2424 21554 2452 21966
rect 2516 21894 2544 23582
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2608 21690 2636 23598
rect 2700 22574 2728 23718
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2792 21554 2820 24550
rect 2884 23497 2912 26726
rect 2976 26353 3004 27270
rect 3056 27056 3108 27062
rect 3056 26998 3108 27004
rect 2962 26344 3018 26353
rect 2962 26279 3018 26288
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2870 23488 2926 23497
rect 2870 23423 2926 23432
rect 2976 23186 3004 26182
rect 3068 25906 3096 26998
rect 3160 26246 3188 29294
rect 3698 29200 3754 30000
rect 4526 29200 4582 30000
rect 5354 29200 5410 30000
rect 6182 29200 6238 30000
rect 7010 29200 7066 30000
rect 7838 29200 7894 30000
rect 8666 29200 8722 30000
rect 9494 29322 9550 30000
rect 10322 29322 10378 30000
rect 9494 29294 9628 29322
rect 9494 29200 9550 29294
rect 3712 27962 3740 29200
rect 3974 28928 4030 28937
rect 3974 28863 4030 28872
rect 3528 27934 3740 27962
rect 3240 27532 3292 27538
rect 3240 27474 3292 27480
rect 3252 26314 3280 27474
rect 3528 26994 3556 27934
rect 3988 27878 4016 28863
rect 4066 28248 4122 28257
rect 4066 28183 4122 28192
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3664 27772 3972 27781
rect 3664 27770 3670 27772
rect 3726 27770 3750 27772
rect 3806 27770 3830 27772
rect 3886 27770 3910 27772
rect 3966 27770 3972 27772
rect 3726 27718 3728 27770
rect 3908 27718 3910 27770
rect 3664 27716 3670 27718
rect 3726 27716 3750 27718
rect 3806 27716 3830 27718
rect 3886 27716 3910 27718
rect 3966 27716 3972 27718
rect 3664 27707 3972 27716
rect 4080 27674 4108 28183
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 27062 4108 27270
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4540 26994 4568 29200
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5368 27418 5396 29200
rect 5724 27464 5776 27470
rect 5170 27024 5226 27033
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 4528 26988 4580 26994
rect 5170 26959 5172 26968
rect 4528 26930 4580 26936
rect 5224 26959 5226 26968
rect 5172 26930 5224 26936
rect 5276 26926 5304 27406
rect 5368 27390 5488 27418
rect 5724 27406 5776 27412
rect 6092 27464 6144 27470
rect 6092 27406 6144 27412
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5368 27130 5396 27270
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5264 26920 5316 26926
rect 4066 26888 4122 26897
rect 5264 26862 5316 26868
rect 4066 26823 4122 26832
rect 3664 26684 3972 26693
rect 3664 26682 3670 26684
rect 3726 26682 3750 26684
rect 3806 26682 3830 26684
rect 3886 26682 3910 26684
rect 3966 26682 3972 26684
rect 3726 26630 3728 26682
rect 3908 26630 3910 26682
rect 3664 26628 3670 26630
rect 3726 26628 3750 26630
rect 3806 26628 3830 26630
rect 3886 26628 3910 26630
rect 3966 26628 3972 26630
rect 3664 26619 3972 26628
rect 4080 26586 4108 26823
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 5368 26353 5396 26726
rect 5460 26382 5488 27390
rect 5736 26382 5764 27406
rect 5448 26376 5500 26382
rect 5354 26344 5410 26353
rect 3240 26308 3292 26314
rect 3240 26250 3292 26256
rect 3332 26308 3384 26314
rect 5448 26318 5500 26324
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5354 26279 5410 26288
rect 3332 26250 3384 26256
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3252 26042 3280 26250
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 3056 25900 3108 25906
rect 3056 25842 3108 25848
rect 3068 25786 3096 25842
rect 3068 25758 3188 25786
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2884 22506 2912 23054
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2884 21962 2912 22442
rect 2872 21956 2924 21962
rect 2872 21898 2924 21904
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2976 20890 3004 22986
rect 3068 22438 3096 25638
rect 3160 23866 3188 25758
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 3160 23118 3188 23462
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 3160 21690 3188 22918
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 3148 21480 3200 21486
rect 3146 21448 3148 21457
rect 3200 21448 3202 21457
rect 3146 21383 3202 21392
rect 3252 21146 3280 25638
rect 3344 24750 3372 26250
rect 4804 26240 4856 26246
rect 4066 26208 4122 26217
rect 4804 26182 4856 26188
rect 4066 26143 4122 26152
rect 4080 25838 4108 26143
rect 4252 25900 4304 25906
rect 4436 25900 4488 25906
rect 4304 25860 4436 25888
rect 4252 25842 4304 25848
rect 4436 25842 4488 25848
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3436 25537 3464 25706
rect 3608 25696 3660 25702
rect 3528 25656 3608 25684
rect 3422 25528 3478 25537
rect 3422 25463 3478 25472
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3344 21010 3372 24686
rect 3436 24138 3464 24822
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3436 23322 3464 24074
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3436 22234 3464 22646
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3528 21536 3556 25656
rect 3608 25638 3660 25644
rect 3664 25596 3972 25605
rect 3664 25594 3670 25596
rect 3726 25594 3750 25596
rect 3806 25594 3830 25596
rect 3886 25594 3910 25596
rect 3966 25594 3972 25596
rect 3726 25542 3728 25594
rect 3908 25542 3910 25594
rect 3664 25540 3670 25542
rect 3726 25540 3750 25542
rect 3806 25540 3830 25542
rect 3886 25540 3910 25542
rect 3966 25540 3972 25542
rect 3664 25531 3972 25540
rect 4264 25430 4292 25842
rect 4252 25424 4304 25430
rect 4252 25366 4304 25372
rect 4528 25424 4580 25430
rect 4528 25366 4580 25372
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 4080 24818 4108 25162
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3620 24614 3648 24754
rect 4264 24698 4292 25230
rect 4080 24670 4292 24698
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3664 24508 3972 24517
rect 3664 24506 3670 24508
rect 3726 24506 3750 24508
rect 3806 24506 3830 24508
rect 3886 24506 3910 24508
rect 3966 24506 3972 24508
rect 3726 24454 3728 24506
rect 3908 24454 3910 24506
rect 3664 24452 3670 24454
rect 3726 24452 3750 24454
rect 3806 24452 3830 24454
rect 3886 24452 3910 24454
rect 3966 24452 3972 24454
rect 3664 24443 3972 24452
rect 3608 24200 3660 24206
rect 4080 24177 4108 24670
rect 4540 24614 4568 25366
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4252 24608 4304 24614
rect 4252 24550 4304 24556
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4172 24206 4200 24550
rect 4264 24410 4292 24550
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4160 24200 4212 24206
rect 3608 24142 3660 24148
rect 4066 24168 4122 24177
rect 3620 23633 3648 24142
rect 4160 24142 4212 24148
rect 4066 24103 4122 24112
rect 4172 23866 4200 24142
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 3606 23624 3662 23633
rect 3606 23559 3662 23568
rect 3664 23420 3972 23429
rect 3664 23418 3670 23420
rect 3726 23418 3750 23420
rect 3806 23418 3830 23420
rect 3886 23418 3910 23420
rect 3966 23418 3972 23420
rect 3726 23366 3728 23418
rect 3908 23366 3910 23418
rect 3664 23364 3670 23366
rect 3726 23364 3750 23366
rect 3806 23364 3830 23366
rect 3886 23364 3910 23366
rect 3966 23364 3972 23366
rect 3664 23355 3972 23364
rect 4080 23050 4108 23802
rect 4356 23225 4384 24550
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4448 24138 4476 24346
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 4158 23216 4214 23225
rect 4158 23151 4214 23160
rect 4342 23216 4398 23225
rect 4342 23151 4398 23160
rect 4172 23118 4200 23151
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 23044 4120 23050
rect 4068 22986 4120 22992
rect 4172 22930 4200 23054
rect 4172 22902 4292 22930
rect 4066 22808 4122 22817
rect 4066 22743 4122 22752
rect 4080 22642 4108 22743
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3882 22536 3938 22545
rect 3882 22471 3884 22480
rect 3936 22471 3938 22480
rect 3884 22442 3936 22448
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 3664 22332 3972 22341
rect 3664 22330 3670 22332
rect 3726 22330 3750 22332
rect 3806 22330 3830 22332
rect 3886 22330 3910 22332
rect 3966 22330 3972 22332
rect 3726 22278 3728 22330
rect 3908 22278 3910 22330
rect 3664 22276 3670 22278
rect 3726 22276 3750 22278
rect 3806 22276 3830 22278
rect 3886 22276 3910 22278
rect 3966 22276 3972 22278
rect 3664 22267 3972 22276
rect 3882 22128 3938 22137
rect 3882 22063 3938 22072
rect 4068 22092 4120 22098
rect 3896 22030 3924 22063
rect 4068 22034 4120 22040
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3436 21508 3556 21536
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 2884 20874 3004 20890
rect 2872 20868 3004 20874
rect 2924 20862 3004 20868
rect 2872 20810 2924 20816
rect 3436 20806 3464 21508
rect 4080 21434 4108 22034
rect 4172 21554 4200 22374
rect 4264 22098 4292 22902
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 4448 21690 4476 23666
rect 4632 23118 4660 25094
rect 4816 24886 4844 26182
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 4724 23798 4752 24210
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 22438 4660 22918
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4080 21406 4200 21434
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 4172 20942 4200 21406
rect 4632 21010 4660 22170
rect 4724 22098 4752 23734
rect 4908 23254 4936 25094
rect 5092 24993 5120 25230
rect 5078 24984 5134 24993
rect 5078 24919 5134 24928
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4896 23248 4948 23254
rect 4802 23216 4858 23225
rect 4896 23190 4948 23196
rect 4802 23151 4858 23160
rect 4816 23050 4844 23151
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 5000 22166 5028 24686
rect 5092 24614 5120 24754
rect 5354 24712 5410 24721
rect 5264 24676 5316 24682
rect 5354 24647 5356 24656
rect 5264 24618 5316 24624
rect 5408 24647 5410 24656
rect 5356 24618 5408 24624
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5276 24562 5304 24618
rect 5276 24534 5396 24562
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 5092 23798 5120 24142
rect 5368 24138 5396 24534
rect 5460 24410 5488 26318
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5172 24064 5224 24070
rect 5170 24032 5172 24041
rect 5224 24032 5226 24041
rect 5170 23967 5226 23976
rect 5368 23798 5396 24074
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5264 23656 5316 23662
rect 5262 23624 5264 23633
rect 5356 23656 5408 23662
rect 5316 23624 5318 23633
rect 5356 23598 5408 23604
rect 5262 23559 5318 23568
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5184 22778 5212 22918
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5276 22556 5304 23559
rect 5368 23526 5396 23598
rect 5460 23594 5488 24210
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5368 23186 5396 23462
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5460 23050 5488 23530
rect 5448 23044 5500 23050
rect 5448 22986 5500 22992
rect 5356 22568 5408 22574
rect 5276 22528 5356 22556
rect 5356 22510 5408 22516
rect 5368 22234 5396 22510
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 4988 22160 5040 22166
rect 4988 22102 5040 22108
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 3424 20800 3476 20806
rect 3054 20768 3110 20777
rect 3424 20742 3476 20748
rect 3054 20703 3110 20712
rect 3068 20466 3096 20703
rect 4816 20602 4844 21966
rect 5368 21690 5396 22170
rect 5460 22137 5488 22986
rect 5446 22128 5502 22137
rect 5446 22063 5502 22072
rect 5552 22094 5580 25978
rect 5632 25220 5684 25226
rect 5632 25162 5684 25168
rect 5644 24206 5672 25162
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5552 22066 5672 22094
rect 5644 22030 5672 22066
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 4908 21146 4936 21626
rect 5828 21418 5856 24006
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5920 23322 5948 23666
rect 6104 23322 6132 27406
rect 6196 25906 6224 29200
rect 6828 27600 6880 27606
rect 7024 27588 7052 29200
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 6880 27560 7052 27588
rect 7194 27568 7250 27577
rect 6828 27542 6880 27548
rect 7194 27503 7250 27512
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6276 27396 6328 27402
rect 6276 27338 6328 27344
rect 6184 25900 6236 25906
rect 6184 25842 6236 25848
rect 6288 25498 6316 27338
rect 6378 27228 6686 27237
rect 6378 27226 6384 27228
rect 6440 27226 6464 27228
rect 6520 27226 6544 27228
rect 6600 27226 6624 27228
rect 6680 27226 6686 27228
rect 6440 27174 6442 27226
rect 6622 27174 6624 27226
rect 6378 27172 6384 27174
rect 6440 27172 6464 27174
rect 6520 27172 6544 27174
rect 6600 27172 6624 27174
rect 6680 27172 6686 27174
rect 6378 27163 6686 27172
rect 6644 26920 6696 26926
rect 6748 26897 6776 27406
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 6840 26994 6868 27338
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6644 26862 6696 26868
rect 6734 26888 6790 26897
rect 6656 26314 6684 26862
rect 6734 26823 6790 26832
rect 6932 26586 6960 27338
rect 7010 27160 7066 27169
rect 7010 27095 7066 27104
rect 7024 27062 7052 27095
rect 7012 27056 7064 27062
rect 7012 26998 7064 27004
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 6736 26580 6788 26586
rect 6920 26580 6972 26586
rect 6788 26540 6868 26568
rect 6736 26522 6788 26528
rect 6734 26480 6790 26489
rect 6840 26466 6868 26540
rect 6920 26522 6972 26528
rect 6840 26438 6960 26466
rect 6734 26415 6790 26424
rect 6748 26382 6776 26415
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6644 26308 6696 26314
rect 6644 26250 6696 26256
rect 6378 26140 6686 26149
rect 6378 26138 6384 26140
rect 6440 26138 6464 26140
rect 6520 26138 6544 26140
rect 6600 26138 6624 26140
rect 6680 26138 6686 26140
rect 6440 26086 6442 26138
rect 6622 26086 6624 26138
rect 6378 26084 6384 26086
rect 6440 26084 6464 26086
rect 6520 26084 6544 26086
rect 6600 26084 6624 26086
rect 6680 26084 6686 26086
rect 6378 26075 6686 26084
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6274 25392 6330 25401
rect 6274 25327 6330 25336
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6196 24138 6224 24890
rect 6288 24818 6316 25327
rect 6932 25294 6960 26438
rect 7024 25906 7052 26726
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6378 25052 6686 25061
rect 6378 25050 6384 25052
rect 6440 25050 6464 25052
rect 6520 25050 6544 25052
rect 6600 25050 6624 25052
rect 6680 25050 6686 25052
rect 6440 24998 6442 25050
rect 6622 24998 6624 25050
rect 6378 24996 6384 24998
rect 6440 24996 6464 24998
rect 6520 24996 6544 24998
rect 6600 24996 6624 24998
rect 6680 24996 6686 24998
rect 6378 24987 6686 24996
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6644 24336 6696 24342
rect 6642 24304 6644 24313
rect 6696 24304 6698 24313
rect 6642 24239 6698 24248
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6196 23866 6224 24074
rect 6378 23964 6686 23973
rect 6378 23962 6384 23964
rect 6440 23962 6464 23964
rect 6520 23962 6544 23964
rect 6600 23962 6624 23964
rect 6680 23962 6686 23964
rect 6440 23910 6442 23962
rect 6622 23910 6624 23962
rect 6378 23908 6384 23910
rect 6440 23908 6464 23910
rect 6520 23908 6544 23910
rect 6600 23908 6624 23910
rect 6680 23908 6686 23910
rect 6378 23899 6686 23908
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6734 23760 6790 23769
rect 6734 23695 6736 23704
rect 6788 23695 6790 23704
rect 6736 23666 6788 23672
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6104 22642 6132 23054
rect 6378 22876 6686 22885
rect 6378 22874 6384 22876
rect 6440 22874 6464 22876
rect 6520 22874 6544 22876
rect 6600 22874 6624 22876
rect 6680 22874 6686 22876
rect 6440 22822 6442 22874
rect 6622 22822 6624 22874
rect 6378 22820 6384 22822
rect 6440 22820 6464 22822
rect 6520 22820 6544 22822
rect 6600 22820 6624 22822
rect 6680 22820 6686 22822
rect 6378 22811 6686 22820
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 6748 22506 6776 23054
rect 6840 22710 6868 23462
rect 6932 23254 6960 25230
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 7116 22778 7144 24822
rect 7208 24342 7236 27503
rect 7286 27024 7342 27033
rect 7286 26959 7342 26968
rect 7196 24336 7248 24342
rect 7196 24278 7248 24284
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6736 22500 6788 22506
rect 6736 22442 6788 22448
rect 7300 22098 7328 26959
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7392 26586 7420 26726
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7484 24818 7512 27814
rect 7564 27668 7616 27674
rect 7564 27610 7616 27616
rect 7576 24818 7604 27610
rect 7656 27056 7708 27062
rect 7656 26998 7708 27004
rect 7748 27056 7800 27062
rect 7852 27033 7880 29200
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8022 27160 8078 27169
rect 8022 27095 8024 27104
rect 8076 27095 8078 27104
rect 8024 27066 8076 27072
rect 8208 27056 8260 27062
rect 7748 26998 7800 27004
rect 7838 27024 7894 27033
rect 7668 26586 7696 26998
rect 7760 26897 7788 26998
rect 8208 26998 8260 27004
rect 7838 26959 7894 26968
rect 7746 26888 7802 26897
rect 7746 26823 7802 26832
rect 8220 26586 8248 26998
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 7748 26512 7800 26518
rect 7748 26454 7800 26460
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7668 25430 7696 25638
rect 7656 25424 7708 25430
rect 7656 25366 7708 25372
rect 7760 25294 7788 26454
rect 8220 26314 8248 26522
rect 8298 26344 8354 26353
rect 8208 26308 8260 26314
rect 8404 26314 8432 27270
rect 8484 26852 8536 26858
rect 8484 26794 8536 26800
rect 8298 26279 8354 26288
rect 8392 26308 8444 26314
rect 8208 26250 8260 26256
rect 7838 25800 7894 25809
rect 7838 25735 7894 25744
rect 7852 25498 7880 25735
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 8312 24818 8340 26279
rect 8392 26250 8444 26256
rect 8496 25294 8524 26794
rect 8680 26450 8708 29200
rect 9092 27772 9400 27781
rect 9092 27770 9098 27772
rect 9154 27770 9178 27772
rect 9234 27770 9258 27772
rect 9314 27770 9338 27772
rect 9394 27770 9400 27772
rect 9154 27718 9156 27770
rect 9336 27718 9338 27770
rect 9092 27716 9098 27718
rect 9154 27716 9178 27718
rect 9234 27716 9258 27718
rect 9314 27716 9338 27718
rect 9394 27716 9400 27718
rect 9092 27707 9400 27716
rect 8944 26852 8996 26858
rect 8944 26794 8996 26800
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8956 26330 8984 26794
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9092 26684 9400 26693
rect 9092 26682 9098 26684
rect 9154 26682 9178 26684
rect 9234 26682 9258 26684
rect 9314 26682 9338 26684
rect 9394 26682 9400 26684
rect 9154 26630 9156 26682
rect 9336 26630 9338 26682
rect 9092 26628 9098 26630
rect 9154 26628 9178 26630
rect 9234 26628 9258 26630
rect 9314 26628 9338 26630
rect 9394 26628 9400 26630
rect 9092 26619 9400 26628
rect 9126 26344 9182 26353
rect 8864 25770 8892 26318
rect 8956 26302 9126 26330
rect 9126 26279 9182 26288
rect 9140 25974 9168 26279
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 8852 25764 8904 25770
rect 8852 25706 8904 25712
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8864 24954 8892 25706
rect 9092 25596 9400 25605
rect 9092 25594 9098 25596
rect 9154 25594 9178 25596
rect 9234 25594 9258 25596
rect 9314 25594 9338 25596
rect 9394 25594 9400 25596
rect 9154 25542 9156 25594
rect 9336 25542 9338 25594
rect 9092 25540 9098 25542
rect 9154 25540 9178 25542
rect 9234 25540 9258 25542
rect 9314 25540 9338 25542
rect 9394 25540 9400 25542
rect 9092 25531 9400 25540
rect 8852 24948 8904 24954
rect 8852 24890 8904 24896
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 7484 24342 7512 24754
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8588 24342 8616 24550
rect 9092 24508 9400 24517
rect 9092 24506 9098 24508
rect 9154 24506 9178 24508
rect 9234 24506 9258 24508
rect 9314 24506 9338 24508
rect 9394 24506 9400 24508
rect 9154 24454 9156 24506
rect 9336 24454 9338 24506
rect 9092 24452 9098 24454
rect 9154 24452 9178 24454
rect 9234 24452 9258 24454
rect 9314 24452 9338 24454
rect 9394 24452 9400 24454
rect 9092 24443 9400 24452
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 9508 24206 9536 26726
rect 9600 24410 9628 29294
rect 9968 29294 10378 29322
rect 9968 27130 9996 29294
rect 10322 29200 10378 29294
rect 11150 29200 11206 30000
rect 11978 29200 12034 30000
rect 12806 29200 12862 30000
rect 13634 29322 13690 30000
rect 13634 29294 13768 29322
rect 13634 29200 13690 29294
rect 10796 27402 11100 27418
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 10784 27396 11112 27402
rect 10836 27390 11060 27396
rect 10784 27338 10836 27344
rect 11060 27338 11112 27344
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10060 27010 10088 27066
rect 9968 26982 10088 27010
rect 9770 26616 9826 26625
rect 9770 26551 9826 26560
rect 9784 26518 9812 26551
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9772 26512 9824 26518
rect 9772 26454 9824 26460
rect 9862 26480 9918 26489
rect 9692 25945 9720 26454
rect 9862 26415 9918 26424
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 9678 25936 9734 25945
rect 9678 25871 9734 25880
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9692 24682 9720 25774
rect 9784 25770 9812 26318
rect 9772 25764 9824 25770
rect 9772 25706 9824 25712
rect 9784 25362 9812 25706
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9876 24682 9904 26415
rect 9968 26246 9996 26982
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 9956 26240 10008 26246
rect 9956 26182 10008 26188
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9968 24614 9996 26182
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 10060 24274 10088 26522
rect 10152 26042 10180 27270
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 10336 25906 10364 27338
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 27112 10732 27270
rect 10704 27084 11008 27112
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10784 26308 10836 26314
rect 10428 26268 10784 26296
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10336 25294 10364 25842
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10428 24410 10456 26268
rect 10784 26250 10836 26256
rect 10506 25936 10562 25945
rect 10506 25871 10508 25880
rect 10560 25871 10562 25880
rect 10508 25842 10560 25848
rect 10612 25214 10824 25242
rect 10612 25158 10640 25214
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 10508 24880 10560 24886
rect 10704 24868 10732 25094
rect 10560 24840 10732 24868
rect 10508 24822 10560 24828
rect 10692 24744 10744 24750
rect 10520 24692 10692 24698
rect 10520 24686 10744 24692
rect 10520 24670 10732 24686
rect 10520 24614 10548 24670
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10692 24608 10744 24614
rect 10796 24562 10824 25214
rect 10744 24556 10824 24562
rect 10692 24550 10824 24556
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 8116 23792 8168 23798
rect 8116 23734 8168 23740
rect 8128 22642 8156 23734
rect 9092 23420 9400 23429
rect 9092 23418 9098 23420
rect 9154 23418 9178 23420
rect 9234 23418 9258 23420
rect 9314 23418 9338 23420
rect 9394 23418 9400 23420
rect 9154 23366 9156 23418
rect 9336 23366 9338 23418
rect 9092 23364 9098 23366
rect 9154 23364 9178 23366
rect 9234 23364 9258 23366
rect 9314 23364 9338 23366
rect 9394 23364 9400 23366
rect 9092 23355 9400 23364
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 9092 22332 9400 22341
rect 9092 22330 9098 22332
rect 9154 22330 9178 22332
rect 9234 22330 9258 22332
rect 9314 22330 9338 22332
rect 9394 22330 9400 22332
rect 9154 22278 9156 22330
rect 9336 22278 9338 22330
rect 9092 22276 9098 22278
rect 9154 22276 9178 22278
rect 9234 22276 9258 22278
rect 9314 22276 9338 22278
rect 9394 22276 9400 22278
rect 9092 22267 9400 22276
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 9876 21554 9904 23258
rect 10520 22094 10548 24550
rect 10704 24534 10824 24550
rect 10888 23866 10916 26930
rect 10980 24954 11008 27084
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 11072 25702 11100 25978
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11072 25226 11100 25638
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11164 24410 11192 29200
rect 11992 27674 12020 29200
rect 11980 27668 12032 27674
rect 11980 27610 12032 27616
rect 12820 27554 12848 29200
rect 12716 27532 12768 27538
rect 12820 27526 13032 27554
rect 12716 27474 12768 27480
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11716 27130 11744 27270
rect 11806 27228 12114 27237
rect 11806 27226 11812 27228
rect 11868 27226 11892 27228
rect 11948 27226 11972 27228
rect 12028 27226 12052 27228
rect 12108 27226 12114 27228
rect 11868 27174 11870 27226
rect 12050 27174 12052 27226
rect 11806 27172 11812 27174
rect 11868 27172 11892 27174
rect 11948 27172 11972 27174
rect 12028 27172 12052 27174
rect 12108 27172 12114 27174
rect 11806 27163 12114 27172
rect 12544 27130 12572 27406
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11428 26920 11480 26926
rect 11242 26888 11298 26897
rect 11428 26862 11480 26868
rect 11242 26823 11298 26832
rect 11256 26790 11284 26823
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11440 26382 11468 26862
rect 11532 26625 11560 26930
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11518 26616 11574 26625
rect 11518 26551 11574 26560
rect 11244 26376 11296 26382
rect 11428 26376 11480 26382
rect 11244 26318 11296 26324
rect 11334 26344 11390 26353
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 11256 23730 11284 26318
rect 11428 26318 11480 26324
rect 11334 26279 11390 26288
rect 11348 24206 11376 26279
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11440 24138 11468 25910
rect 11532 25158 11560 26551
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11624 24818 11652 26726
rect 11992 26518 12020 26998
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 11980 26512 12032 26518
rect 11978 26480 11980 26489
rect 12164 26512 12216 26518
rect 12032 26480 12034 26489
rect 11704 26444 11756 26450
rect 12164 26454 12216 26460
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 11978 26415 12034 26424
rect 11704 26386 11756 26392
rect 11716 26042 11744 26386
rect 11992 26228 12020 26415
rect 12176 26382 12204 26454
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 11992 26200 12204 26228
rect 11806 26140 12114 26149
rect 11806 26138 11812 26140
rect 11868 26138 11892 26140
rect 11948 26138 11972 26140
rect 12028 26138 12052 26140
rect 12108 26138 12114 26140
rect 11868 26086 11870 26138
rect 12050 26086 12052 26138
rect 11806 26084 11812 26086
rect 11868 26084 11892 26086
rect 11948 26084 11972 26086
rect 12028 26084 12052 26086
rect 12108 26084 12114 26086
rect 11806 26075 12114 26084
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 12176 25974 12204 26200
rect 12268 26042 12296 26318
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 11808 25498 11836 25638
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 12268 25294 12296 25638
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 11806 25052 12114 25061
rect 11806 25050 11812 25052
rect 11868 25050 11892 25052
rect 11948 25050 11972 25052
rect 12028 25050 12052 25052
rect 12108 25050 12114 25052
rect 11868 24998 11870 25050
rect 12050 24998 12052 25050
rect 11806 24996 11812 24998
rect 11868 24996 11892 24998
rect 11948 24996 11972 24998
rect 12028 24996 12052 24998
rect 12108 24996 12114 24998
rect 11806 24987 12114 24996
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12360 24274 12388 26454
rect 12452 25702 12480 26726
rect 12728 26432 12756 27474
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12912 26790 12940 27406
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12636 26404 12756 26432
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12544 25294 12572 26182
rect 12636 25294 12664 26404
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12728 25430 12756 26250
rect 12716 25424 12768 25430
rect 12716 25366 12768 25372
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12820 24818 12848 26522
rect 12912 25809 12940 26726
rect 13004 26382 13032 27526
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13096 27062 13124 27406
rect 13176 27396 13228 27402
rect 13176 27338 13228 27344
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 13188 26994 13216 27338
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 13096 26518 13124 26862
rect 13084 26512 13136 26518
rect 13084 26454 13136 26460
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 12898 25800 12954 25809
rect 12898 25735 12954 25744
rect 13082 25800 13138 25809
rect 13082 25735 13138 25744
rect 13096 25702 13124 25735
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 13188 24342 13216 26250
rect 13280 25906 13308 27406
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13280 25498 13308 25842
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13372 25294 13400 26182
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13464 25226 13492 27270
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13556 25702 13584 26318
rect 13648 26314 13676 26998
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13740 25786 13768 29294
rect 14462 29200 14518 30000
rect 15290 29200 15346 30000
rect 16118 29322 16174 30000
rect 16118 29294 16528 29322
rect 16118 29200 16174 29294
rect 14476 27962 14504 29200
rect 14384 27934 14504 27962
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 14016 26994 14044 27542
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13832 26450 13860 26930
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13924 26042 13952 26726
rect 14200 26489 14228 27474
rect 14384 26518 14412 27934
rect 14520 27772 14828 27781
rect 14520 27770 14526 27772
rect 14582 27770 14606 27772
rect 14662 27770 14686 27772
rect 14742 27770 14766 27772
rect 14822 27770 14828 27772
rect 14582 27718 14584 27770
rect 14764 27718 14766 27770
rect 14520 27716 14526 27718
rect 14582 27716 14606 27718
rect 14662 27716 14686 27718
rect 14742 27716 14766 27718
rect 14822 27716 14828 27718
rect 14520 27707 14828 27716
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14476 26772 14504 27610
rect 14648 27532 14700 27538
rect 14568 27492 14648 27520
rect 14568 27130 14596 27492
rect 14648 27474 14700 27480
rect 14648 27396 14700 27402
rect 14648 27338 14700 27344
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14660 26790 14688 27338
rect 14924 26852 14976 26858
rect 14924 26794 14976 26800
rect 14444 26744 14504 26772
rect 14648 26784 14700 26790
rect 14444 26586 14472 26744
rect 14648 26726 14700 26732
rect 14520 26684 14828 26693
rect 14520 26682 14526 26684
rect 14582 26682 14606 26684
rect 14662 26682 14686 26684
rect 14742 26682 14766 26684
rect 14822 26682 14828 26684
rect 14582 26630 14584 26682
rect 14764 26630 14766 26682
rect 14520 26628 14526 26630
rect 14582 26628 14606 26630
rect 14662 26628 14686 26630
rect 14742 26628 14766 26630
rect 14822 26628 14828 26630
rect 14520 26619 14828 26628
rect 14444 26580 14516 26586
rect 14444 26540 14464 26580
rect 14464 26522 14516 26528
rect 14280 26512 14332 26518
rect 14186 26480 14242 26489
rect 14280 26454 14332 26460
rect 14372 26512 14424 26518
rect 14372 26454 14424 26460
rect 14186 26415 14242 26424
rect 14200 26314 14228 26415
rect 14292 26353 14320 26454
rect 14278 26344 14334 26353
rect 14188 26308 14240 26314
rect 14278 26279 14334 26288
rect 14188 26250 14240 26256
rect 14280 26240 14332 26246
rect 14280 26182 14332 26188
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13912 25832 13964 25838
rect 13740 25780 13912 25786
rect 13740 25774 13964 25780
rect 13740 25758 13952 25774
rect 14292 25770 14320 26182
rect 14372 25900 14424 25906
rect 14476 25888 14504 26522
rect 14936 26314 14964 26794
rect 15304 26382 15332 29200
rect 15752 27396 15804 27402
rect 15752 27338 15804 27344
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 15764 26246 15792 27338
rect 16500 26976 16528 29294
rect 16946 29200 17002 30000
rect 17774 29200 17830 30000
rect 18602 29200 18658 30000
rect 19430 29200 19486 30000
rect 20258 29200 20314 30000
rect 21086 29200 21142 30000
rect 21914 29200 21970 30000
rect 22742 29322 22798 30000
rect 22480 29294 22798 29322
rect 16960 27606 16988 29200
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 17040 27464 17092 27470
rect 17788 27452 17816 29200
rect 18616 27470 18644 29200
rect 19444 27606 19472 29200
rect 20272 27962 20300 29200
rect 20272 27934 20392 27962
rect 19948 27772 20256 27781
rect 19948 27770 19954 27772
rect 20010 27770 20034 27772
rect 20090 27770 20114 27772
rect 20170 27770 20194 27772
rect 20250 27770 20256 27772
rect 20010 27718 20012 27770
rect 20192 27718 20194 27770
rect 19948 27716 19954 27718
rect 20010 27716 20034 27718
rect 20090 27716 20114 27718
rect 20170 27716 20194 27718
rect 20250 27716 20256 27718
rect 19948 27707 20256 27716
rect 20364 27606 20392 27934
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 20352 27600 20404 27606
rect 20352 27542 20404 27548
rect 17960 27464 18012 27470
rect 17788 27424 17960 27452
rect 17040 27406 17092 27412
rect 17960 27406 18012 27412
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 16580 26988 16632 26994
rect 16500 26948 16580 26976
rect 16580 26930 16632 26936
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 25974 15792 26182
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 14424 25860 14504 25888
rect 14372 25842 14424 25848
rect 14384 25809 14412 25842
rect 14370 25800 14426 25809
rect 14280 25764 14332 25770
rect 14370 25735 14426 25744
rect 14280 25706 14332 25712
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 14292 24886 14320 25706
rect 14520 25596 14828 25605
rect 14520 25594 14526 25596
rect 14582 25594 14606 25596
rect 14662 25594 14686 25596
rect 14742 25594 14766 25596
rect 14822 25594 14828 25596
rect 14582 25542 14584 25594
rect 14764 25542 14766 25594
rect 14520 25540 14526 25542
rect 14582 25540 14606 25542
rect 14662 25540 14686 25542
rect 14742 25540 14766 25542
rect 14822 25540 14828 25542
rect 14520 25531 14828 25540
rect 14280 24880 14332 24886
rect 14280 24822 14332 24828
rect 17052 24750 17080 27406
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 17234 27228 17542 27237
rect 17234 27226 17240 27228
rect 17296 27226 17320 27228
rect 17376 27226 17400 27228
rect 17456 27226 17480 27228
rect 17536 27226 17542 27228
rect 17296 27174 17298 27226
rect 17478 27174 17480 27226
rect 17234 27172 17240 27174
rect 17296 27172 17320 27174
rect 17376 27172 17400 27174
rect 17456 27172 17480 27174
rect 17536 27172 17542 27174
rect 17234 27163 17542 27172
rect 18156 27062 18184 27270
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 20364 26994 20392 27542
rect 20536 27464 20588 27470
rect 20536 27406 20588 27412
rect 20548 27130 20576 27406
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 18144 26920 18196 26926
rect 20536 26920 20588 26926
rect 18144 26862 18196 26868
rect 20534 26888 20536 26897
rect 20588 26888 20590 26897
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17972 26450 18000 26726
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 18156 26314 18184 26862
rect 21100 26858 21128 29200
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 20534 26823 20590 26832
rect 21088 26852 21140 26858
rect 21088 26794 21140 26800
rect 19948 26684 20256 26693
rect 19948 26682 19954 26684
rect 20010 26682 20034 26684
rect 20090 26682 20114 26684
rect 20170 26682 20194 26684
rect 20250 26682 20256 26684
rect 20010 26630 20012 26682
rect 20192 26630 20194 26682
rect 19948 26628 19954 26630
rect 20010 26628 20034 26630
rect 20090 26628 20114 26630
rect 20170 26628 20194 26630
rect 20250 26628 20256 26630
rect 19948 26619 20256 26628
rect 19432 26376 19484 26382
rect 19430 26344 19432 26353
rect 20628 26376 20680 26382
rect 19484 26344 19486 26353
rect 18144 26308 18196 26314
rect 20628 26318 20680 26324
rect 19430 26279 19486 26288
rect 18144 26250 18196 26256
rect 17234 26140 17542 26149
rect 17234 26138 17240 26140
rect 17296 26138 17320 26140
rect 17376 26138 17400 26140
rect 17456 26138 17480 26140
rect 17536 26138 17542 26140
rect 17296 26086 17298 26138
rect 17478 26086 17480 26138
rect 17234 26084 17240 26086
rect 17296 26084 17320 26086
rect 17376 26084 17400 26086
rect 17456 26084 17480 26086
rect 17536 26084 17542 26086
rect 17234 26075 17542 26084
rect 18156 26042 18184 26250
rect 19524 26240 19576 26246
rect 19524 26182 19576 26188
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19444 25809 19472 25842
rect 19430 25800 19486 25809
rect 19430 25735 19486 25744
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17234 25052 17542 25061
rect 17234 25050 17240 25052
rect 17296 25050 17320 25052
rect 17376 25050 17400 25052
rect 17456 25050 17480 25052
rect 17536 25050 17542 25052
rect 17296 24998 17298 25050
rect 17478 24998 17480 25050
rect 17234 24996 17240 24998
rect 17296 24996 17320 24998
rect 17376 24996 17400 24998
rect 17456 24996 17480 24998
rect 17536 24996 17542 24998
rect 17234 24987 17542 24996
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 14520 24508 14828 24517
rect 14520 24506 14526 24508
rect 14582 24506 14606 24508
rect 14662 24506 14686 24508
rect 14742 24506 14766 24508
rect 14822 24506 14828 24508
rect 14582 24454 14584 24506
rect 14764 24454 14766 24506
rect 14520 24452 14526 24454
rect 14582 24452 14606 24454
rect 14662 24452 14686 24454
rect 14742 24452 14766 24454
rect 14822 24452 14828 24454
rect 14520 24443 14828 24452
rect 17420 24410 17448 24754
rect 17788 24614 17816 25094
rect 19352 24886 19380 25434
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11428 24132 11480 24138
rect 11428 24074 11480 24080
rect 11806 23964 12114 23973
rect 11806 23962 11812 23964
rect 11868 23962 11892 23964
rect 11948 23962 11972 23964
rect 12028 23962 12052 23964
rect 12108 23962 12114 23964
rect 11868 23910 11870 23962
rect 12050 23910 12052 23962
rect 11806 23908 11812 23910
rect 11868 23908 11892 23910
rect 11948 23908 11972 23910
rect 12028 23908 12052 23910
rect 12108 23908 12114 23910
rect 11806 23899 12114 23908
rect 12360 23798 12388 24210
rect 17234 23964 17542 23973
rect 17234 23962 17240 23964
rect 17296 23962 17320 23964
rect 17376 23962 17400 23964
rect 17456 23962 17480 23964
rect 17536 23962 17542 23964
rect 17296 23910 17298 23962
rect 17478 23910 17480 23962
rect 17234 23908 17240 23910
rect 17296 23908 17320 23910
rect 17376 23908 17400 23910
rect 17456 23908 17480 23910
rect 17536 23908 17542 23910
rect 17234 23899 17542 23908
rect 17604 23866 17632 24346
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 16672 23792 16724 23798
rect 16672 23734 16724 23740
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 14520 23420 14828 23429
rect 14520 23418 14526 23420
rect 14582 23418 14606 23420
rect 14662 23418 14686 23420
rect 14742 23418 14766 23420
rect 14822 23418 14828 23420
rect 14582 23366 14584 23418
rect 14764 23366 14766 23418
rect 14520 23364 14526 23366
rect 14582 23364 14606 23366
rect 14662 23364 14686 23366
rect 14742 23364 14766 23366
rect 14822 23364 14828 23366
rect 14520 23355 14828 23364
rect 16684 23050 16712 23734
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 11806 22876 12114 22885
rect 11806 22874 11812 22876
rect 11868 22874 11892 22876
rect 11948 22874 11972 22876
rect 12028 22874 12052 22876
rect 12108 22874 12114 22876
rect 11868 22822 11870 22874
rect 12050 22822 12052 22874
rect 11806 22820 11812 22822
rect 11868 22820 11892 22822
rect 11948 22820 11972 22822
rect 12028 22820 12052 22822
rect 12108 22820 12114 22822
rect 11806 22811 12114 22820
rect 14520 22332 14828 22341
rect 14520 22330 14526 22332
rect 14582 22330 14606 22332
rect 14662 22330 14686 22332
rect 14742 22330 14766 22332
rect 14822 22330 14828 22332
rect 14582 22278 14584 22330
rect 14764 22278 14766 22330
rect 14520 22276 14526 22278
rect 14582 22276 14606 22278
rect 14662 22276 14686 22278
rect 14742 22276 14766 22278
rect 14822 22276 14828 22278
rect 14520 22267 14828 22276
rect 16868 22166 16896 23258
rect 17040 23248 17092 23254
rect 17038 23216 17040 23225
rect 17092 23216 17094 23225
rect 17038 23151 17094 23160
rect 17236 23050 17264 23666
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17696 22982 17724 24142
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17234 22876 17542 22885
rect 17234 22874 17240 22876
rect 17296 22874 17320 22876
rect 17376 22874 17400 22876
rect 17456 22874 17480 22876
rect 17536 22874 17542 22876
rect 17296 22822 17298 22874
rect 17478 22822 17480 22874
rect 17234 22820 17240 22822
rect 17296 22820 17320 22822
rect 17376 22820 17400 22822
rect 17456 22820 17480 22822
rect 17536 22820 17542 22822
rect 17234 22811 17542 22820
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 16856 22160 16908 22166
rect 17604 22137 17632 22374
rect 16856 22102 16908 22108
rect 17590 22128 17646 22137
rect 10600 22094 10652 22098
rect 10520 22092 10652 22094
rect 10520 22066 10600 22092
rect 10600 22034 10652 22040
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 10336 21010 10364 21286
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 7116 20534 7144 20742
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7392 20466 7420 20946
rect 10428 20942 10456 21830
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 20097 2452 20198
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 2410 20088 2466 20097
rect 3664 20091 3972 20100
rect 2410 20023 2466 20032
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 1504 18737 1532 19790
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17218 1532 17614
rect 1596 17377 1624 19110
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1582 17368 1638 17377
rect 1582 17303 1638 17312
rect 1504 17190 1624 17218
rect 1596 17134 1624 17190
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16794 1624 17070
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15162 1624 15438
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1688 12442 1716 17546
rect 1872 16590 1900 19450
rect 2240 19417 2268 19790
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 2226 19408 2282 19417
rect 2226 19343 2282 19352
rect 2410 19408 2466 19417
rect 2410 19343 2412 19352
rect 2464 19343 2466 19352
rect 2412 19314 2464 19320
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2792 18766 2820 19110
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 1950 18184 2006 18193
rect 1950 18119 2006 18128
rect 2044 18148 2096 18154
rect 1964 18086 1992 18119
rect 2044 18090 2096 18096
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1780 13530 1808 15370
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 14074 1992 15302
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2056 13734 2084 18090
rect 2240 16590 2268 18294
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 15366 2268 16526
rect 2332 15366 2360 18158
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 16250 2636 17614
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2424 13530 2452 15438
rect 2608 15094 2636 16186
rect 2700 15609 2728 17478
rect 2792 16697 2820 18702
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2778 16688 2834 16697
rect 2778 16623 2834 16632
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2608 14906 2636 15030
rect 2608 14878 2728 14906
rect 2596 14816 2648 14822
rect 2516 14764 2596 14770
rect 2516 14758 2648 14764
rect 2516 14742 2636 14758
rect 2516 13870 2544 14742
rect 2700 14634 2728 14878
rect 2608 14606 2728 14634
rect 2608 13938 2636 14606
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1780 11354 1808 13466
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1964 12374 1992 13262
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12714 2360 13194
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12850 2452 13126
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 2226 11928 2282 11937
rect 2516 11898 2544 13806
rect 2608 12714 2636 13874
rect 2700 13530 2728 14214
rect 2792 13802 2820 15642
rect 2884 14414 2912 18566
rect 3068 18290 3096 18906
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3344 18426 3372 18702
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2976 17338 3004 18226
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2976 17066 3004 17274
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2976 16114 3004 16730
rect 3068 16454 3096 18226
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2976 15570 3004 16050
rect 3054 15600 3110 15609
rect 2964 15564 3016 15570
rect 3054 15535 3110 15544
rect 2964 15506 3016 15512
rect 3068 15502 3096 15535
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2976 14074 3004 15370
rect 3054 15328 3110 15337
rect 3054 15263 3110 15272
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2884 13394 2912 13670
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2792 12442 2820 13223
rect 2884 12850 2912 13330
rect 3068 12850 3096 15263
rect 3160 14074 3188 17070
rect 3252 15706 3280 17546
rect 3344 16250 3372 18158
rect 3436 17202 3464 19654
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 3516 18080 3568 18086
rect 3514 18048 3516 18057
rect 3568 18048 3570 18057
rect 3514 17983 3570 17992
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3252 15314 3280 15506
rect 3344 15434 3372 16186
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3252 15286 3372 15314
rect 3344 14958 3372 15286
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3330 14784 3386 14793
rect 3330 14719 3386 14728
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3160 13190 3188 13738
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12918 3188 13126
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2226 11863 2282 11872
rect 2504 11892 2556 11898
rect 2240 11762 2268 11863
rect 2504 11834 2556 11840
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 9178 1532 11086
rect 2792 10810 2820 12174
rect 3160 11830 3188 12582
rect 3252 12306 3280 14486
rect 3344 13938 3372 14719
rect 3436 14346 3464 16594
rect 3528 15162 3556 17138
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 4080 15502 4108 16934
rect 4172 16017 4200 17002
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4158 16008 4214 16017
rect 4158 15943 4214 15952
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15570 4200 15846
rect 4264 15638 4292 16934
rect 4356 16794 4384 17478
rect 4448 17270 4476 17478
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16454 4384 16526
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4342 15600 4398 15609
rect 4160 15564 4212 15570
rect 4632 15570 4660 18634
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 15706 4752 17138
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16658 4936 16934
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4816 15638 4844 16390
rect 4908 16046 4936 16594
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4342 15535 4398 15544
rect 4620 15564 4672 15570
rect 4160 15506 4212 15512
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 14952 3568 14958
rect 3620 14929 3648 15302
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3516 14894 3568 14900
rect 3606 14920 3662 14929
rect 3528 14498 3556 14894
rect 3606 14855 3662 14864
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3528 14482 3740 14498
rect 3528 14476 3752 14482
rect 3528 14470 3700 14476
rect 3700 14418 3752 14424
rect 3884 14408 3936 14414
rect 3514 14376 3570 14385
rect 3424 14340 3476 14346
rect 3884 14350 3936 14356
rect 3514 14311 3570 14320
rect 3424 14282 3476 14288
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3344 13530 3372 13874
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3436 12782 3464 14282
rect 3528 13326 3556 14311
rect 3896 13977 3924 14350
rect 3988 14074 4016 14554
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3882 13968 3938 13977
rect 3792 13932 3844 13938
rect 3882 13903 3938 13912
rect 3792 13874 3844 13880
rect 3804 13734 3832 13874
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3528 12617 3556 12786
rect 3514 12608 3570 12617
rect 3514 12543 3570 12552
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 4080 12442 4108 14962
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14346 4200 14894
rect 4356 14600 4384 15535
rect 4620 15506 4672 15512
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4264 14572 4384 14600
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4264 13938 4292 14572
rect 4342 14512 4398 14521
rect 4342 14447 4344 14456
rect 4396 14447 4398 14456
rect 4344 14418 4396 14424
rect 4540 14074 4568 15438
rect 4816 14890 4844 15574
rect 5000 15162 5028 17614
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5184 16522 5212 17274
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5078 15736 5134 15745
rect 5078 15671 5080 15680
rect 5132 15671 5134 15680
rect 5080 15642 5132 15648
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5184 15026 5212 16458
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 15706 5304 16390
rect 5552 16046 5580 16526
rect 5736 16046 5764 18838
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 5816 17604 5868 17610
rect 5816 17546 5868 17552
rect 5828 16454 5856 17546
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 6378 17371 6686 17380
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6012 16590 6040 16730
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6012 16250 6040 16390
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5552 15026 5580 15846
rect 5920 15706 5948 16118
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6104 15502 6132 16662
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6196 15366 6224 16118
rect 6288 15570 6316 16390
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 15706 6592 16050
rect 6748 15910 6776 18770
rect 7392 18714 7420 20402
rect 8772 20262 8800 20878
rect 10612 20330 10640 21490
rect 11716 21146 11744 21966
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 11716 19514 11744 21082
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 12544 19378 12572 20198
rect 13372 19378 13400 20402
rect 16868 20398 16896 22102
rect 17590 22063 17646 22072
rect 17696 21962 17724 22918
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17788 21894 17816 24550
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23798 17908 24006
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 18064 23730 18092 24686
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17880 22574 17908 23190
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18248 22778 18276 23122
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 17788 21350 17816 21830
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17788 21010 17816 21286
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 17788 20262 17816 20946
rect 18340 20806 18368 22986
rect 18616 22030 18644 23462
rect 18708 22642 18736 24550
rect 19352 24426 19380 24822
rect 19260 24398 19380 24426
rect 19444 24410 19472 25230
rect 19432 24404 19484 24410
rect 19260 24206 19288 24398
rect 19432 24346 19484 24352
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19248 24200 19300 24206
rect 19352 24177 19380 24210
rect 19248 24142 19300 24148
rect 19338 24168 19394 24177
rect 19076 23730 19104 24142
rect 19338 24103 19394 24112
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19352 23730 19380 23802
rect 19430 23760 19486 23769
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 19340 23724 19392 23730
rect 19536 23730 19564 26182
rect 19708 25900 19760 25906
rect 19708 25842 19760 25848
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19628 24410 19656 24550
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19430 23695 19486 23704
rect 19524 23724 19576 23730
rect 19340 23666 19392 23672
rect 19076 23050 19104 23666
rect 19444 23594 19472 23695
rect 19524 23666 19576 23672
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19444 22964 19472 23258
rect 19628 23118 19656 24142
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19306 22936 19472 22964
rect 19524 22976 19576 22982
rect 19522 22944 19524 22953
rect 19576 22944 19578 22953
rect 19306 22778 19334 22936
rect 19522 22879 19578 22888
rect 19720 22778 19748 25842
rect 19892 25832 19944 25838
rect 19812 25792 19892 25820
rect 19812 25498 19840 25792
rect 19892 25774 19944 25780
rect 19948 25596 20256 25605
rect 19948 25594 19954 25596
rect 20010 25594 20034 25596
rect 20090 25594 20114 25596
rect 20170 25594 20194 25596
rect 20250 25594 20256 25596
rect 20010 25542 20012 25594
rect 20192 25542 20194 25594
rect 19948 25540 19954 25542
rect 20010 25540 20034 25542
rect 20090 25540 20114 25542
rect 20170 25540 20194 25542
rect 20250 25540 20256 25542
rect 19948 25531 20256 25540
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 20076 25152 20128 25158
rect 20128 25100 20208 25106
rect 20076 25094 20208 25100
rect 20088 25078 20208 25094
rect 20180 24886 20208 25078
rect 20168 24880 20220 24886
rect 20168 24822 20220 24828
rect 19800 24676 19852 24682
rect 19800 24618 19852 24624
rect 19812 23633 19840 24618
rect 19948 24508 20256 24517
rect 19948 24506 19954 24508
rect 20010 24506 20034 24508
rect 20090 24506 20114 24508
rect 20170 24506 20194 24508
rect 20250 24506 20256 24508
rect 20010 24454 20012 24506
rect 20192 24454 20194 24506
rect 19948 24452 19954 24454
rect 20010 24452 20034 24454
rect 20090 24452 20114 24454
rect 20170 24452 20194 24454
rect 20250 24452 20256 24454
rect 19948 24443 20256 24452
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19996 24070 20024 24142
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19798 23624 19854 23633
rect 19798 23559 19854 23568
rect 19996 23508 20024 24006
rect 19812 23480 20024 23508
rect 19812 22982 19840 23480
rect 19948 23420 20256 23429
rect 19948 23418 19954 23420
rect 20010 23418 20034 23420
rect 20090 23418 20114 23420
rect 20170 23418 20194 23420
rect 20250 23418 20256 23420
rect 20010 23366 20012 23418
rect 20192 23366 20194 23418
rect 19948 23364 19954 23366
rect 20010 23364 20034 23366
rect 20090 23364 20114 23366
rect 20170 23364 20194 23366
rect 20250 23364 20256 23366
rect 19948 23355 20256 23364
rect 20364 23322 20392 25842
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20444 25492 20496 25498
rect 20444 25434 20496 25440
rect 20456 23866 20484 25434
rect 20548 25294 20576 25638
rect 20536 25288 20588 25294
rect 20640 25265 20668 26318
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20904 26308 20956 26314
rect 20904 26250 20956 26256
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20536 25230 20588 25236
rect 20626 25256 20682 25265
rect 20626 25191 20682 25200
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 19294 22772 19346 22778
rect 19294 22714 19346 22720
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19432 22704 19484 22710
rect 19430 22672 19432 22681
rect 19484 22672 19486 22681
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 19248 22636 19300 22642
rect 19430 22607 19486 22616
rect 19248 22578 19300 22584
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18892 22030 18920 22374
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21690 18828 21830
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 19260 21350 19288 22578
rect 19904 22488 19932 23054
rect 20088 22778 20116 23122
rect 20456 23118 20484 23462
rect 20444 23112 20496 23118
rect 20350 23080 20406 23089
rect 20444 23054 20496 23060
rect 20350 23015 20406 23024
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 19812 22460 19932 22488
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19706 22400 19762 22409
rect 19340 22160 19392 22166
rect 19392 22120 19472 22148
rect 19340 22102 19392 22108
rect 19340 22024 19392 22030
rect 19338 21992 19340 22001
rect 19392 21992 19394 22001
rect 19338 21927 19394 21936
rect 19444 21622 19472 22120
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19432 21480 19484 21486
rect 19430 21448 19432 21457
rect 19524 21480 19576 21486
rect 19484 21448 19486 21457
rect 19524 21422 19576 21428
rect 19430 21383 19486 21392
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19536 21146 19564 21422
rect 19628 21418 19656 22374
rect 19706 22335 19762 22344
rect 19616 21412 19668 21418
rect 19616 21354 19668 21360
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19720 20942 19748 22335
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19812 20874 19840 22460
rect 20088 22438 20116 22714
rect 20180 22642 20208 22714
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19948 22332 20256 22341
rect 19948 22330 19954 22332
rect 20010 22330 20034 22332
rect 20090 22330 20114 22332
rect 20170 22330 20194 22332
rect 20250 22330 20256 22332
rect 20010 22278 20012 22330
rect 20192 22278 20194 22330
rect 19948 22276 19954 22278
rect 20010 22276 20034 22278
rect 20090 22276 20114 22278
rect 20170 22276 20194 22278
rect 20250 22276 20256 22278
rect 19948 22267 20256 22276
rect 19892 22024 19944 22030
rect 19890 21992 19892 22001
rect 19944 21992 19946 22001
rect 19890 21927 19946 21936
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19996 21486 20024 21898
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 21622 20300 21830
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 14292 20058 14320 20198
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 19628 19922 19656 20742
rect 20364 20466 20392 23015
rect 20548 22817 20576 25094
rect 20640 23186 20668 25094
rect 20732 24410 20760 25366
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20534 22808 20590 22817
rect 20732 22794 20760 23802
rect 20534 22743 20590 22752
rect 20640 22766 20760 22794
rect 20442 21992 20498 22001
rect 20442 21927 20498 21936
rect 20456 20466 20484 21927
rect 20548 21894 20576 22743
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20548 20534 20576 21558
rect 20640 21146 20668 22766
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20732 21962 20760 22646
rect 20824 22234 20852 26250
rect 20916 25498 20944 26250
rect 21088 25832 21140 25838
rect 21088 25774 21140 25780
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 21100 24954 21128 25774
rect 21284 25702 21312 26250
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21088 24948 21140 24954
rect 21088 24890 21140 24896
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20916 23050 20944 23258
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20902 22128 20958 22137
rect 20902 22063 20958 22072
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20732 21486 20760 21558
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 20824 20058 20852 21490
rect 20916 20602 20944 22063
rect 21008 20942 21036 24822
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21100 22166 21128 23122
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 21192 22030 21220 25638
rect 21284 24342 21312 25638
rect 21272 24336 21324 24342
rect 21272 24278 21324 24284
rect 21376 23730 21404 27270
rect 21456 26784 21508 26790
rect 21456 26726 21508 26732
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21468 24721 21496 26726
rect 21560 24818 21588 26726
rect 21638 26480 21694 26489
rect 21638 26415 21640 26424
rect 21692 26415 21694 26424
rect 21640 26386 21692 26392
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 25226 21680 26250
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21640 25220 21692 25226
rect 21640 25162 21692 25168
rect 21640 24948 21692 24954
rect 21640 24890 21692 24896
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21454 24712 21510 24721
rect 21454 24647 21510 24656
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21284 23118 21312 23462
rect 21376 23186 21404 23666
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21362 22944 21418 22953
rect 21284 22098 21312 22918
rect 21362 22879 21418 22888
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 21622 21128 21830
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 21284 21554 21312 21626
rect 21272 21548 21324 21554
rect 21376 21536 21404 22879
rect 21468 22710 21496 24550
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21560 22574 21588 23598
rect 21652 22778 21680 24890
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21560 21962 21588 22510
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21456 21548 21508 21554
rect 21376 21508 21456 21536
rect 21272 21490 21324 21496
rect 21456 21490 21508 21496
rect 21560 21146 21588 21898
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21362 20904 21418 20913
rect 21362 20839 21418 20848
rect 21270 20632 21326 20641
rect 20904 20596 20956 20602
rect 21270 20567 21326 20576
rect 20904 20538 20956 20544
rect 21284 20262 21312 20567
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 21376 19854 21404 20839
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 12394 19372 12446 19378
rect 12268 19332 12394 19360
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 9508 18766 9536 19246
rect 12268 19174 12296 19332
rect 12394 19314 12446 19320
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 9496 18760 9548 18766
rect 7392 18686 7512 18714
rect 9496 18702 9548 18708
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18358 7420 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7484 18290 7512 18686
rect 9508 18426 9536 18702
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 16998 7512 18226
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6748 15638 6776 15846
rect 6736 15632 6788 15638
rect 6932 15609 6960 16118
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 6736 15574 6788 15580
rect 6918 15600 6974 15609
rect 6276 15564 6328 15570
rect 6918 15535 6974 15544
rect 6276 15506 6328 15512
rect 10980 15502 11008 19110
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 21560 18970 21588 21082
rect 21652 20874 21680 22714
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 21744 20602 21772 25842
rect 21836 23769 21864 27270
rect 21928 27062 21956 29200
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21928 24410 21956 26250
rect 22112 25770 22140 27406
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 21822 23760 21878 23769
rect 21822 23695 21878 23704
rect 21836 22642 21864 23695
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21928 22438 21956 24346
rect 22020 24206 22048 25638
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22112 23254 22140 24754
rect 22204 24138 22232 26930
rect 22480 26042 22508 29294
rect 22742 29200 22798 29294
rect 22662 27228 22970 27237
rect 22662 27226 22668 27228
rect 22724 27226 22748 27228
rect 22804 27226 22828 27228
rect 22884 27226 22908 27228
rect 22964 27226 22970 27228
rect 22724 27174 22726 27226
rect 22906 27174 22908 27226
rect 22662 27172 22668 27174
rect 22724 27172 22748 27174
rect 22804 27172 22828 27174
rect 22884 27172 22908 27174
rect 22964 27172 22970 27174
rect 22662 27163 22970 27172
rect 22662 26140 22970 26149
rect 22662 26138 22668 26140
rect 22724 26138 22748 26140
rect 22804 26138 22828 26140
rect 22884 26138 22908 26140
rect 22964 26138 22970 26140
rect 22724 26086 22726 26138
rect 22906 26086 22908 26138
rect 22662 26084 22668 26086
rect 22724 26084 22748 26086
rect 22804 26084 22828 26086
rect 22884 26084 22908 26086
rect 22964 26084 22970 26086
rect 22662 26075 22970 26084
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22388 24750 22416 25230
rect 22662 25052 22970 25061
rect 22662 25050 22668 25052
rect 22724 25050 22748 25052
rect 22804 25050 22828 25052
rect 22884 25050 22908 25052
rect 22964 25050 22970 25052
rect 22724 24998 22726 25050
rect 22906 24998 22908 25050
rect 22662 24996 22668 24998
rect 22724 24996 22748 24998
rect 22804 24996 22828 24998
rect 22884 24996 22908 24998
rect 22964 24996 22970 24998
rect 22662 24987 22970 24996
rect 22376 24744 22428 24750
rect 22376 24686 22428 24692
rect 22388 24206 22416 24686
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22100 23248 22152 23254
rect 22204 23225 22232 23666
rect 22388 23662 22416 24142
rect 22662 23964 22970 23973
rect 22662 23962 22668 23964
rect 22724 23962 22748 23964
rect 22804 23962 22828 23964
rect 22884 23962 22908 23964
rect 22964 23962 22970 23964
rect 22724 23910 22726 23962
rect 22906 23910 22908 23962
rect 22662 23908 22668 23910
rect 22724 23908 22748 23910
rect 22804 23908 22828 23910
rect 22884 23908 22908 23910
rect 22964 23908 22970 23910
rect 22662 23899 22970 23908
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22100 23190 22152 23196
rect 22190 23216 22246 23225
rect 22190 23151 22246 23160
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21928 20058 21956 22374
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22020 20369 22048 21286
rect 22006 20360 22062 20369
rect 22006 20295 22062 20304
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22020 19281 22048 19314
rect 22006 19272 22062 19281
rect 22006 19207 22062 19216
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22020 16561 22048 16594
rect 22006 16552 22062 16561
rect 22006 16487 22062 16496
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 22112 16250 22140 22578
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22204 20058 22232 21558
rect 22296 21146 22324 23054
rect 22662 22876 22970 22885
rect 22662 22874 22668 22876
rect 22724 22874 22748 22876
rect 22804 22874 22828 22876
rect 22884 22874 22908 22876
rect 22964 22874 22970 22876
rect 22724 22822 22726 22874
rect 22906 22822 22908 22874
rect 22662 22820 22668 22822
rect 22724 22820 22748 22822
rect 22804 22820 22828 22822
rect 22884 22820 22908 22822
rect 22964 22820 22970 22822
rect 22662 22811 22970 22820
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22296 19825 22324 20198
rect 22282 19816 22338 19825
rect 22282 19751 22338 19760
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 17882 22232 19110
rect 22284 18760 22336 18766
rect 22282 18728 22284 18737
rect 22336 18728 22338 18737
rect 22282 18663 22338 18672
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 22282 18184 22338 18193
rect 22282 18119 22284 18128
rect 22336 18119 22338 18128
rect 22284 18090 22336 18096
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22284 17672 22336 17678
rect 22282 17640 22284 17649
rect 22336 17640 22338 17649
rect 22282 17575 22338 17584
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 22282 17096 22338 17105
rect 22282 17031 22284 17040
rect 22336 17031 22338 17040
rect 22284 17002 22336 17008
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22112 16017 22140 16050
rect 22098 16008 22154 16017
rect 22098 15943 22154 15952
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 10968 15496 11020 15502
rect 22284 15496 22336 15502
rect 10968 15438 11020 15444
rect 22282 15464 22284 15473
rect 22336 15464 22338 15473
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14346 4844 14826
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4448 13530 4476 13874
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4632 12986 4660 14214
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 6748 13870 6776 15438
rect 22282 15399 22338 15408
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 6378 11931 6686 11940
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 11257 2912 11494
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 2870 11248 2926 11257
rect 2870 11183 2926 11192
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10577 1624 10610
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9897 1624 9998
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 1582 9208 1638 9217
rect 3664 9211 3972 9220
rect 1492 9172 1544 9178
rect 1582 9143 1638 9152
rect 1492 9114 1544 9120
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1780 8537 1808 8910
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 1766 8528 1822 8537
rect 1766 8463 1822 8472
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 1584 7880 1636 7886
rect 1582 7848 1584 7857
rect 1636 7848 1638 7857
rect 1582 7783 1638 7792
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 7484 6322 7512 15302
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 22282 14920 22338 14929
rect 22282 14855 22284 14864
rect 22336 14855 22338 14864
rect 22284 14826 22336 14832
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 22284 13864 22336 13870
rect 22282 13832 22284 13841
rect 22336 13832 22338 13841
rect 22282 13767 22338 13776
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 22284 13320 22336 13326
rect 22282 13288 22284 13297
rect 22336 13288 22338 13297
rect 22282 13223 22338 13232
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 22284 12232 22336 12238
rect 22282 12200 22284 12209
rect 22336 12200 22338 12209
rect 22282 12135 22338 12144
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 22282 11656 22338 11665
rect 22282 11591 22284 11600
rect 22336 11591 22338 11600
rect 22284 11562 22336 11568
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 22282 10568 22338 10577
rect 22282 10503 22284 10512
rect 22336 10503 22338 10512
rect 22284 10474 22336 10480
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 22284 10056 22336 10062
rect 22282 10024 22284 10033
rect 22336 10024 22338 10033
rect 22282 9959 22338 9968
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 22284 8968 22336 8974
rect 22282 8936 22284 8945
rect 22336 8936 22338 8945
rect 22282 8871 22338 8880
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 22282 8392 22338 8401
rect 22282 8327 22284 8336
rect 22336 8327 22338 8336
rect 22284 8298 22336 8304
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 22282 7304 22338 7313
rect 22282 7239 22284 7248
rect 22336 7239 22338 7248
rect 22284 7210 22336 7216
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 22284 6792 22336 6798
rect 22282 6760 22284 6769
rect 22336 6760 22338 6769
rect 22282 6695 22338 6704
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5817 1716 6054
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 22284 5704 22336 5710
rect 22282 5672 22284 5681
rect 22336 5672 22338 5681
rect 22282 5607 22338 5616
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 1584 5160 1636 5166
rect 1582 5128 1584 5137
rect 1636 5128 1638 5137
rect 1582 5063 1638 5072
rect 22282 5128 22338 5137
rect 22282 5063 22284 5072
rect 22336 5063 22338 5072
rect 22284 5034 22336 5040
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 22282 4040 22338 4049
rect 22282 3975 22284 3984
rect 22336 3975 22338 3984
rect 22284 3946 22336 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3777 1624 3878
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 1582 3768 1638 3777
rect 3664 3771 3972 3780
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 1582 3703 1638 3712
rect 1584 3528 1636 3534
rect 22284 3528 22336 3534
rect 1584 3470 1636 3476
rect 22282 3496 22284 3505
rect 22336 3496 22338 3505
rect 1596 3097 1624 3470
rect 22282 3431 22338 3440
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 1057 1440 2790
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1596 1737 1624 2382
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
rect 1582 1728 1638 1737
rect 1582 1663 1638 1672
rect 1398 1048 1454 1057
rect 1398 983 1454 992
<< via2 >>
rect 1214 25336 1270 25392
rect 2502 24792 2558 24848
rect 2686 24656 2742 24712
rect 2686 24248 2742 24304
rect 2594 23976 2650 24032
rect 2134 21684 2190 21720
rect 2134 21664 2136 21684
rect 2136 21664 2188 21684
rect 2188 21664 2190 21684
rect 2962 26288 3018 26344
rect 2870 23432 2926 23488
rect 3974 28872 4030 28928
rect 4066 28192 4122 28248
rect 3670 27770 3726 27772
rect 3750 27770 3806 27772
rect 3830 27770 3886 27772
rect 3910 27770 3966 27772
rect 3670 27718 3716 27770
rect 3716 27718 3726 27770
rect 3750 27718 3780 27770
rect 3780 27718 3792 27770
rect 3792 27718 3806 27770
rect 3830 27718 3844 27770
rect 3844 27718 3856 27770
rect 3856 27718 3886 27770
rect 3910 27718 3920 27770
rect 3920 27718 3966 27770
rect 3670 27716 3726 27718
rect 3750 27716 3806 27718
rect 3830 27716 3886 27718
rect 3910 27716 3966 27718
rect 5170 26988 5226 27024
rect 5170 26968 5172 26988
rect 5172 26968 5224 26988
rect 5224 26968 5226 26988
rect 4066 26832 4122 26888
rect 3670 26682 3726 26684
rect 3750 26682 3806 26684
rect 3830 26682 3886 26684
rect 3910 26682 3966 26684
rect 3670 26630 3716 26682
rect 3716 26630 3726 26682
rect 3750 26630 3780 26682
rect 3780 26630 3792 26682
rect 3792 26630 3806 26682
rect 3830 26630 3844 26682
rect 3844 26630 3856 26682
rect 3856 26630 3886 26682
rect 3910 26630 3920 26682
rect 3920 26630 3966 26682
rect 3670 26628 3726 26630
rect 3750 26628 3806 26630
rect 3830 26628 3886 26630
rect 3910 26628 3966 26630
rect 5354 26288 5410 26344
rect 3146 21428 3148 21448
rect 3148 21428 3200 21448
rect 3200 21428 3202 21448
rect 3146 21392 3202 21428
rect 4066 26152 4122 26208
rect 3422 25472 3478 25528
rect 3670 25594 3726 25596
rect 3750 25594 3806 25596
rect 3830 25594 3886 25596
rect 3910 25594 3966 25596
rect 3670 25542 3716 25594
rect 3716 25542 3726 25594
rect 3750 25542 3780 25594
rect 3780 25542 3792 25594
rect 3792 25542 3806 25594
rect 3830 25542 3844 25594
rect 3844 25542 3856 25594
rect 3856 25542 3886 25594
rect 3910 25542 3920 25594
rect 3920 25542 3966 25594
rect 3670 25540 3726 25542
rect 3750 25540 3806 25542
rect 3830 25540 3886 25542
rect 3910 25540 3966 25542
rect 3670 24506 3726 24508
rect 3750 24506 3806 24508
rect 3830 24506 3886 24508
rect 3910 24506 3966 24508
rect 3670 24454 3716 24506
rect 3716 24454 3726 24506
rect 3750 24454 3780 24506
rect 3780 24454 3792 24506
rect 3792 24454 3806 24506
rect 3830 24454 3844 24506
rect 3844 24454 3856 24506
rect 3856 24454 3886 24506
rect 3910 24454 3920 24506
rect 3920 24454 3966 24506
rect 3670 24452 3726 24454
rect 3750 24452 3806 24454
rect 3830 24452 3886 24454
rect 3910 24452 3966 24454
rect 4066 24112 4122 24168
rect 3606 23568 3662 23624
rect 3670 23418 3726 23420
rect 3750 23418 3806 23420
rect 3830 23418 3886 23420
rect 3910 23418 3966 23420
rect 3670 23366 3716 23418
rect 3716 23366 3726 23418
rect 3750 23366 3780 23418
rect 3780 23366 3792 23418
rect 3792 23366 3806 23418
rect 3830 23366 3844 23418
rect 3844 23366 3856 23418
rect 3856 23366 3886 23418
rect 3910 23366 3920 23418
rect 3920 23366 3966 23418
rect 3670 23364 3726 23366
rect 3750 23364 3806 23366
rect 3830 23364 3886 23366
rect 3910 23364 3966 23366
rect 4158 23160 4214 23216
rect 4342 23160 4398 23216
rect 4066 22752 4122 22808
rect 3882 22500 3938 22536
rect 3882 22480 3884 22500
rect 3884 22480 3936 22500
rect 3936 22480 3938 22500
rect 3670 22330 3726 22332
rect 3750 22330 3806 22332
rect 3830 22330 3886 22332
rect 3910 22330 3966 22332
rect 3670 22278 3716 22330
rect 3716 22278 3726 22330
rect 3750 22278 3780 22330
rect 3780 22278 3792 22330
rect 3792 22278 3806 22330
rect 3830 22278 3844 22330
rect 3844 22278 3856 22330
rect 3856 22278 3886 22330
rect 3910 22278 3920 22330
rect 3920 22278 3966 22330
rect 3670 22276 3726 22278
rect 3750 22276 3806 22278
rect 3830 22276 3886 22278
rect 3910 22276 3966 22278
rect 3882 22072 3938 22128
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 5078 24928 5134 24984
rect 4802 23160 4858 23216
rect 5354 24676 5410 24712
rect 5354 24656 5356 24676
rect 5356 24656 5408 24676
rect 5408 24656 5410 24676
rect 5170 24012 5172 24032
rect 5172 24012 5224 24032
rect 5224 24012 5226 24032
rect 5170 23976 5226 24012
rect 5262 23604 5264 23624
rect 5264 23604 5316 23624
rect 5316 23604 5318 23624
rect 5262 23568 5318 23604
rect 3054 20712 3110 20768
rect 5446 22072 5502 22128
rect 7194 27512 7250 27568
rect 6384 27226 6440 27228
rect 6464 27226 6520 27228
rect 6544 27226 6600 27228
rect 6624 27226 6680 27228
rect 6384 27174 6430 27226
rect 6430 27174 6440 27226
rect 6464 27174 6494 27226
rect 6494 27174 6506 27226
rect 6506 27174 6520 27226
rect 6544 27174 6558 27226
rect 6558 27174 6570 27226
rect 6570 27174 6600 27226
rect 6624 27174 6634 27226
rect 6634 27174 6680 27226
rect 6384 27172 6440 27174
rect 6464 27172 6520 27174
rect 6544 27172 6600 27174
rect 6624 27172 6680 27174
rect 6734 26832 6790 26888
rect 7010 27104 7066 27160
rect 6734 26424 6790 26480
rect 6384 26138 6440 26140
rect 6464 26138 6520 26140
rect 6544 26138 6600 26140
rect 6624 26138 6680 26140
rect 6384 26086 6430 26138
rect 6430 26086 6440 26138
rect 6464 26086 6494 26138
rect 6494 26086 6506 26138
rect 6506 26086 6520 26138
rect 6544 26086 6558 26138
rect 6558 26086 6570 26138
rect 6570 26086 6600 26138
rect 6624 26086 6634 26138
rect 6634 26086 6680 26138
rect 6384 26084 6440 26086
rect 6464 26084 6520 26086
rect 6544 26084 6600 26086
rect 6624 26084 6680 26086
rect 6274 25336 6330 25392
rect 6384 25050 6440 25052
rect 6464 25050 6520 25052
rect 6544 25050 6600 25052
rect 6624 25050 6680 25052
rect 6384 24998 6430 25050
rect 6430 24998 6440 25050
rect 6464 24998 6494 25050
rect 6494 24998 6506 25050
rect 6506 24998 6520 25050
rect 6544 24998 6558 25050
rect 6558 24998 6570 25050
rect 6570 24998 6600 25050
rect 6624 24998 6634 25050
rect 6634 24998 6680 25050
rect 6384 24996 6440 24998
rect 6464 24996 6520 24998
rect 6544 24996 6600 24998
rect 6624 24996 6680 24998
rect 6642 24284 6644 24304
rect 6644 24284 6696 24304
rect 6696 24284 6698 24304
rect 6642 24248 6698 24284
rect 6384 23962 6440 23964
rect 6464 23962 6520 23964
rect 6544 23962 6600 23964
rect 6624 23962 6680 23964
rect 6384 23910 6430 23962
rect 6430 23910 6440 23962
rect 6464 23910 6494 23962
rect 6494 23910 6506 23962
rect 6506 23910 6520 23962
rect 6544 23910 6558 23962
rect 6558 23910 6570 23962
rect 6570 23910 6600 23962
rect 6624 23910 6634 23962
rect 6634 23910 6680 23962
rect 6384 23908 6440 23910
rect 6464 23908 6520 23910
rect 6544 23908 6600 23910
rect 6624 23908 6680 23910
rect 6734 23724 6790 23760
rect 6734 23704 6736 23724
rect 6736 23704 6788 23724
rect 6788 23704 6790 23724
rect 6384 22874 6440 22876
rect 6464 22874 6520 22876
rect 6544 22874 6600 22876
rect 6624 22874 6680 22876
rect 6384 22822 6430 22874
rect 6430 22822 6440 22874
rect 6464 22822 6494 22874
rect 6494 22822 6506 22874
rect 6506 22822 6520 22874
rect 6544 22822 6558 22874
rect 6558 22822 6570 22874
rect 6570 22822 6600 22874
rect 6624 22822 6634 22874
rect 6634 22822 6680 22874
rect 6384 22820 6440 22822
rect 6464 22820 6520 22822
rect 6544 22820 6600 22822
rect 6624 22820 6680 22822
rect 7286 26968 7342 27024
rect 8022 27124 8078 27160
rect 8022 27104 8024 27124
rect 8024 27104 8076 27124
rect 8076 27104 8078 27124
rect 7838 26968 7894 27024
rect 7746 26832 7802 26888
rect 8298 26288 8354 26344
rect 7838 25744 7894 25800
rect 9098 27770 9154 27772
rect 9178 27770 9234 27772
rect 9258 27770 9314 27772
rect 9338 27770 9394 27772
rect 9098 27718 9144 27770
rect 9144 27718 9154 27770
rect 9178 27718 9208 27770
rect 9208 27718 9220 27770
rect 9220 27718 9234 27770
rect 9258 27718 9272 27770
rect 9272 27718 9284 27770
rect 9284 27718 9314 27770
rect 9338 27718 9348 27770
rect 9348 27718 9394 27770
rect 9098 27716 9154 27718
rect 9178 27716 9234 27718
rect 9258 27716 9314 27718
rect 9338 27716 9394 27718
rect 9098 26682 9154 26684
rect 9178 26682 9234 26684
rect 9258 26682 9314 26684
rect 9338 26682 9394 26684
rect 9098 26630 9144 26682
rect 9144 26630 9154 26682
rect 9178 26630 9208 26682
rect 9208 26630 9220 26682
rect 9220 26630 9234 26682
rect 9258 26630 9272 26682
rect 9272 26630 9284 26682
rect 9284 26630 9314 26682
rect 9338 26630 9348 26682
rect 9348 26630 9394 26682
rect 9098 26628 9154 26630
rect 9178 26628 9234 26630
rect 9258 26628 9314 26630
rect 9338 26628 9394 26630
rect 9126 26288 9182 26344
rect 9098 25594 9154 25596
rect 9178 25594 9234 25596
rect 9258 25594 9314 25596
rect 9338 25594 9394 25596
rect 9098 25542 9144 25594
rect 9144 25542 9154 25594
rect 9178 25542 9208 25594
rect 9208 25542 9220 25594
rect 9220 25542 9234 25594
rect 9258 25542 9272 25594
rect 9272 25542 9284 25594
rect 9284 25542 9314 25594
rect 9338 25542 9348 25594
rect 9348 25542 9394 25594
rect 9098 25540 9154 25542
rect 9178 25540 9234 25542
rect 9258 25540 9314 25542
rect 9338 25540 9394 25542
rect 9098 24506 9154 24508
rect 9178 24506 9234 24508
rect 9258 24506 9314 24508
rect 9338 24506 9394 24508
rect 9098 24454 9144 24506
rect 9144 24454 9154 24506
rect 9178 24454 9208 24506
rect 9208 24454 9220 24506
rect 9220 24454 9234 24506
rect 9258 24454 9272 24506
rect 9272 24454 9284 24506
rect 9284 24454 9314 24506
rect 9338 24454 9348 24506
rect 9348 24454 9394 24506
rect 9098 24452 9154 24454
rect 9178 24452 9234 24454
rect 9258 24452 9314 24454
rect 9338 24452 9394 24454
rect 9770 26560 9826 26616
rect 9862 26424 9918 26480
rect 9678 25880 9734 25936
rect 10506 25900 10562 25936
rect 10506 25880 10508 25900
rect 10508 25880 10560 25900
rect 10560 25880 10562 25900
rect 9098 23418 9154 23420
rect 9178 23418 9234 23420
rect 9258 23418 9314 23420
rect 9338 23418 9394 23420
rect 9098 23366 9144 23418
rect 9144 23366 9154 23418
rect 9178 23366 9208 23418
rect 9208 23366 9220 23418
rect 9220 23366 9234 23418
rect 9258 23366 9272 23418
rect 9272 23366 9284 23418
rect 9284 23366 9314 23418
rect 9338 23366 9348 23418
rect 9348 23366 9394 23418
rect 9098 23364 9154 23366
rect 9178 23364 9234 23366
rect 9258 23364 9314 23366
rect 9338 23364 9394 23366
rect 9098 22330 9154 22332
rect 9178 22330 9234 22332
rect 9258 22330 9314 22332
rect 9338 22330 9394 22332
rect 9098 22278 9144 22330
rect 9144 22278 9154 22330
rect 9178 22278 9208 22330
rect 9208 22278 9220 22330
rect 9220 22278 9234 22330
rect 9258 22278 9272 22330
rect 9272 22278 9284 22330
rect 9284 22278 9314 22330
rect 9338 22278 9348 22330
rect 9348 22278 9394 22330
rect 9098 22276 9154 22278
rect 9178 22276 9234 22278
rect 9258 22276 9314 22278
rect 9338 22276 9394 22278
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 27226 11868 27228
rect 11892 27226 11948 27228
rect 11972 27226 12028 27228
rect 12052 27226 12108 27228
rect 11812 27174 11858 27226
rect 11858 27174 11868 27226
rect 11892 27174 11922 27226
rect 11922 27174 11934 27226
rect 11934 27174 11948 27226
rect 11972 27174 11986 27226
rect 11986 27174 11998 27226
rect 11998 27174 12028 27226
rect 12052 27174 12062 27226
rect 12062 27174 12108 27226
rect 11812 27172 11868 27174
rect 11892 27172 11948 27174
rect 11972 27172 12028 27174
rect 12052 27172 12108 27174
rect 11242 26832 11298 26888
rect 11518 26560 11574 26616
rect 11334 26288 11390 26344
rect 11978 26460 11980 26480
rect 11980 26460 12032 26480
rect 12032 26460 12034 26480
rect 11978 26424 12034 26460
rect 11812 26138 11868 26140
rect 11892 26138 11948 26140
rect 11972 26138 12028 26140
rect 12052 26138 12108 26140
rect 11812 26086 11858 26138
rect 11858 26086 11868 26138
rect 11892 26086 11922 26138
rect 11922 26086 11934 26138
rect 11934 26086 11948 26138
rect 11972 26086 11986 26138
rect 11986 26086 11998 26138
rect 11998 26086 12028 26138
rect 12052 26086 12062 26138
rect 12062 26086 12108 26138
rect 11812 26084 11868 26086
rect 11892 26084 11948 26086
rect 11972 26084 12028 26086
rect 12052 26084 12108 26086
rect 11812 25050 11868 25052
rect 11892 25050 11948 25052
rect 11972 25050 12028 25052
rect 12052 25050 12108 25052
rect 11812 24998 11858 25050
rect 11858 24998 11868 25050
rect 11892 24998 11922 25050
rect 11922 24998 11934 25050
rect 11934 24998 11948 25050
rect 11972 24998 11986 25050
rect 11986 24998 11998 25050
rect 11998 24998 12028 25050
rect 12052 24998 12062 25050
rect 12062 24998 12108 25050
rect 11812 24996 11868 24998
rect 11892 24996 11948 24998
rect 11972 24996 12028 24998
rect 12052 24996 12108 24998
rect 12898 25744 12954 25800
rect 13082 25744 13138 25800
rect 14526 27770 14582 27772
rect 14606 27770 14662 27772
rect 14686 27770 14742 27772
rect 14766 27770 14822 27772
rect 14526 27718 14572 27770
rect 14572 27718 14582 27770
rect 14606 27718 14636 27770
rect 14636 27718 14648 27770
rect 14648 27718 14662 27770
rect 14686 27718 14700 27770
rect 14700 27718 14712 27770
rect 14712 27718 14742 27770
rect 14766 27718 14776 27770
rect 14776 27718 14822 27770
rect 14526 27716 14582 27718
rect 14606 27716 14662 27718
rect 14686 27716 14742 27718
rect 14766 27716 14822 27718
rect 14526 26682 14582 26684
rect 14606 26682 14662 26684
rect 14686 26682 14742 26684
rect 14766 26682 14822 26684
rect 14526 26630 14572 26682
rect 14572 26630 14582 26682
rect 14606 26630 14636 26682
rect 14636 26630 14648 26682
rect 14648 26630 14662 26682
rect 14686 26630 14700 26682
rect 14700 26630 14712 26682
rect 14712 26630 14742 26682
rect 14766 26630 14776 26682
rect 14776 26630 14822 26682
rect 14526 26628 14582 26630
rect 14606 26628 14662 26630
rect 14686 26628 14742 26630
rect 14766 26628 14822 26630
rect 14186 26424 14242 26480
rect 14278 26288 14334 26344
rect 19954 27770 20010 27772
rect 20034 27770 20090 27772
rect 20114 27770 20170 27772
rect 20194 27770 20250 27772
rect 19954 27718 20000 27770
rect 20000 27718 20010 27770
rect 20034 27718 20064 27770
rect 20064 27718 20076 27770
rect 20076 27718 20090 27770
rect 20114 27718 20128 27770
rect 20128 27718 20140 27770
rect 20140 27718 20170 27770
rect 20194 27718 20204 27770
rect 20204 27718 20250 27770
rect 19954 27716 20010 27718
rect 20034 27716 20090 27718
rect 20114 27716 20170 27718
rect 20194 27716 20250 27718
rect 14370 25744 14426 25800
rect 14526 25594 14582 25596
rect 14606 25594 14662 25596
rect 14686 25594 14742 25596
rect 14766 25594 14822 25596
rect 14526 25542 14572 25594
rect 14572 25542 14582 25594
rect 14606 25542 14636 25594
rect 14636 25542 14648 25594
rect 14648 25542 14662 25594
rect 14686 25542 14700 25594
rect 14700 25542 14712 25594
rect 14712 25542 14742 25594
rect 14766 25542 14776 25594
rect 14776 25542 14822 25594
rect 14526 25540 14582 25542
rect 14606 25540 14662 25542
rect 14686 25540 14742 25542
rect 14766 25540 14822 25542
rect 17240 27226 17296 27228
rect 17320 27226 17376 27228
rect 17400 27226 17456 27228
rect 17480 27226 17536 27228
rect 17240 27174 17286 27226
rect 17286 27174 17296 27226
rect 17320 27174 17350 27226
rect 17350 27174 17362 27226
rect 17362 27174 17376 27226
rect 17400 27174 17414 27226
rect 17414 27174 17426 27226
rect 17426 27174 17456 27226
rect 17480 27174 17490 27226
rect 17490 27174 17536 27226
rect 17240 27172 17296 27174
rect 17320 27172 17376 27174
rect 17400 27172 17456 27174
rect 17480 27172 17536 27174
rect 20534 26868 20536 26888
rect 20536 26868 20588 26888
rect 20588 26868 20590 26888
rect 20534 26832 20590 26868
rect 19954 26682 20010 26684
rect 20034 26682 20090 26684
rect 20114 26682 20170 26684
rect 20194 26682 20250 26684
rect 19954 26630 20000 26682
rect 20000 26630 20010 26682
rect 20034 26630 20064 26682
rect 20064 26630 20076 26682
rect 20076 26630 20090 26682
rect 20114 26630 20128 26682
rect 20128 26630 20140 26682
rect 20140 26630 20170 26682
rect 20194 26630 20204 26682
rect 20204 26630 20250 26682
rect 19954 26628 20010 26630
rect 20034 26628 20090 26630
rect 20114 26628 20170 26630
rect 20194 26628 20250 26630
rect 19430 26324 19432 26344
rect 19432 26324 19484 26344
rect 19484 26324 19486 26344
rect 19430 26288 19486 26324
rect 17240 26138 17296 26140
rect 17320 26138 17376 26140
rect 17400 26138 17456 26140
rect 17480 26138 17536 26140
rect 17240 26086 17286 26138
rect 17286 26086 17296 26138
rect 17320 26086 17350 26138
rect 17350 26086 17362 26138
rect 17362 26086 17376 26138
rect 17400 26086 17414 26138
rect 17414 26086 17426 26138
rect 17426 26086 17456 26138
rect 17480 26086 17490 26138
rect 17490 26086 17536 26138
rect 17240 26084 17296 26086
rect 17320 26084 17376 26086
rect 17400 26084 17456 26086
rect 17480 26084 17536 26086
rect 19430 25744 19486 25800
rect 17240 25050 17296 25052
rect 17320 25050 17376 25052
rect 17400 25050 17456 25052
rect 17480 25050 17536 25052
rect 17240 24998 17286 25050
rect 17286 24998 17296 25050
rect 17320 24998 17350 25050
rect 17350 24998 17362 25050
rect 17362 24998 17376 25050
rect 17400 24998 17414 25050
rect 17414 24998 17426 25050
rect 17426 24998 17456 25050
rect 17480 24998 17490 25050
rect 17490 24998 17536 25050
rect 17240 24996 17296 24998
rect 17320 24996 17376 24998
rect 17400 24996 17456 24998
rect 17480 24996 17536 24998
rect 14526 24506 14582 24508
rect 14606 24506 14662 24508
rect 14686 24506 14742 24508
rect 14766 24506 14822 24508
rect 14526 24454 14572 24506
rect 14572 24454 14582 24506
rect 14606 24454 14636 24506
rect 14636 24454 14648 24506
rect 14648 24454 14662 24506
rect 14686 24454 14700 24506
rect 14700 24454 14712 24506
rect 14712 24454 14742 24506
rect 14766 24454 14776 24506
rect 14776 24454 14822 24506
rect 14526 24452 14582 24454
rect 14606 24452 14662 24454
rect 14686 24452 14742 24454
rect 14766 24452 14822 24454
rect 11812 23962 11868 23964
rect 11892 23962 11948 23964
rect 11972 23962 12028 23964
rect 12052 23962 12108 23964
rect 11812 23910 11858 23962
rect 11858 23910 11868 23962
rect 11892 23910 11922 23962
rect 11922 23910 11934 23962
rect 11934 23910 11948 23962
rect 11972 23910 11986 23962
rect 11986 23910 11998 23962
rect 11998 23910 12028 23962
rect 12052 23910 12062 23962
rect 12062 23910 12108 23962
rect 11812 23908 11868 23910
rect 11892 23908 11948 23910
rect 11972 23908 12028 23910
rect 12052 23908 12108 23910
rect 17240 23962 17296 23964
rect 17320 23962 17376 23964
rect 17400 23962 17456 23964
rect 17480 23962 17536 23964
rect 17240 23910 17286 23962
rect 17286 23910 17296 23962
rect 17320 23910 17350 23962
rect 17350 23910 17362 23962
rect 17362 23910 17376 23962
rect 17400 23910 17414 23962
rect 17414 23910 17426 23962
rect 17426 23910 17456 23962
rect 17480 23910 17490 23962
rect 17490 23910 17536 23962
rect 17240 23908 17296 23910
rect 17320 23908 17376 23910
rect 17400 23908 17456 23910
rect 17480 23908 17536 23910
rect 14526 23418 14582 23420
rect 14606 23418 14662 23420
rect 14686 23418 14742 23420
rect 14766 23418 14822 23420
rect 14526 23366 14572 23418
rect 14572 23366 14582 23418
rect 14606 23366 14636 23418
rect 14636 23366 14648 23418
rect 14648 23366 14662 23418
rect 14686 23366 14700 23418
rect 14700 23366 14712 23418
rect 14712 23366 14742 23418
rect 14766 23366 14776 23418
rect 14776 23366 14822 23418
rect 14526 23364 14582 23366
rect 14606 23364 14662 23366
rect 14686 23364 14742 23366
rect 14766 23364 14822 23366
rect 11812 22874 11868 22876
rect 11892 22874 11948 22876
rect 11972 22874 12028 22876
rect 12052 22874 12108 22876
rect 11812 22822 11858 22874
rect 11858 22822 11868 22874
rect 11892 22822 11922 22874
rect 11922 22822 11934 22874
rect 11934 22822 11948 22874
rect 11972 22822 11986 22874
rect 11986 22822 11998 22874
rect 11998 22822 12028 22874
rect 12052 22822 12062 22874
rect 12062 22822 12108 22874
rect 11812 22820 11868 22822
rect 11892 22820 11948 22822
rect 11972 22820 12028 22822
rect 12052 22820 12108 22822
rect 14526 22330 14582 22332
rect 14606 22330 14662 22332
rect 14686 22330 14742 22332
rect 14766 22330 14822 22332
rect 14526 22278 14572 22330
rect 14572 22278 14582 22330
rect 14606 22278 14636 22330
rect 14636 22278 14648 22330
rect 14648 22278 14662 22330
rect 14686 22278 14700 22330
rect 14700 22278 14712 22330
rect 14712 22278 14742 22330
rect 14766 22278 14776 22330
rect 14776 22278 14822 22330
rect 14526 22276 14582 22278
rect 14606 22276 14662 22278
rect 14686 22276 14742 22278
rect 14766 22276 14822 22278
rect 17038 23196 17040 23216
rect 17040 23196 17092 23216
rect 17092 23196 17094 23216
rect 17038 23160 17094 23196
rect 17240 22874 17296 22876
rect 17320 22874 17376 22876
rect 17400 22874 17456 22876
rect 17480 22874 17536 22876
rect 17240 22822 17286 22874
rect 17286 22822 17296 22874
rect 17320 22822 17350 22874
rect 17350 22822 17362 22874
rect 17362 22822 17376 22874
rect 17400 22822 17414 22874
rect 17414 22822 17426 22874
rect 17426 22822 17456 22874
rect 17480 22822 17490 22874
rect 17490 22822 17536 22874
rect 17240 22820 17296 22822
rect 17320 22820 17376 22822
rect 17400 22820 17456 22822
rect 17480 22820 17536 22822
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 2410 20032 2466 20088
rect 1490 18672 1546 18728
rect 1582 17312 1638 17368
rect 2226 19352 2282 19408
rect 2410 19372 2466 19408
rect 2410 19352 2412 19372
rect 2412 19352 2464 19372
rect 2464 19352 2466 19372
rect 1950 18128 2006 18184
rect 2778 16632 2834 16688
rect 2686 15544 2742 15600
rect 2226 11872 2282 11928
rect 3054 15544 3110 15600
rect 3054 15272 3110 15328
rect 2778 13232 2834 13288
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 3514 18028 3516 18048
rect 3516 18028 3568 18048
rect 3568 18028 3570 18048
rect 3514 17992 3570 18028
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 3330 14728 3386 14784
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 4158 15952 4214 16008
rect 4342 15544 4398 15600
rect 3606 14864 3662 14920
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 3514 14320 3570 14376
rect 3882 13912 3938 13968
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3514 12552 3570 12608
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 4342 14476 4398 14512
rect 4342 14456 4344 14476
rect 4344 14456 4396 14476
rect 4396 14456 4398 14476
rect 5078 15700 5134 15736
rect 5078 15680 5080 15700
rect 5080 15680 5132 15700
rect 5132 15680 5134 15700
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 17590 22072 17646 22128
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 19338 24112 19394 24168
rect 19430 23704 19486 23760
rect 19522 22924 19524 22944
rect 19524 22924 19576 22944
rect 19576 22924 19578 22944
rect 19522 22888 19578 22924
rect 19954 25594 20010 25596
rect 20034 25594 20090 25596
rect 20114 25594 20170 25596
rect 20194 25594 20250 25596
rect 19954 25542 20000 25594
rect 20000 25542 20010 25594
rect 20034 25542 20064 25594
rect 20064 25542 20076 25594
rect 20076 25542 20090 25594
rect 20114 25542 20128 25594
rect 20128 25542 20140 25594
rect 20140 25542 20170 25594
rect 20194 25542 20204 25594
rect 20204 25542 20250 25594
rect 19954 25540 20010 25542
rect 20034 25540 20090 25542
rect 20114 25540 20170 25542
rect 20194 25540 20250 25542
rect 19954 24506 20010 24508
rect 20034 24506 20090 24508
rect 20114 24506 20170 24508
rect 20194 24506 20250 24508
rect 19954 24454 20000 24506
rect 20000 24454 20010 24506
rect 20034 24454 20064 24506
rect 20064 24454 20076 24506
rect 20076 24454 20090 24506
rect 20114 24454 20128 24506
rect 20128 24454 20140 24506
rect 20140 24454 20170 24506
rect 20194 24454 20204 24506
rect 20204 24454 20250 24506
rect 19954 24452 20010 24454
rect 20034 24452 20090 24454
rect 20114 24452 20170 24454
rect 20194 24452 20250 24454
rect 19798 23568 19854 23624
rect 19954 23418 20010 23420
rect 20034 23418 20090 23420
rect 20114 23418 20170 23420
rect 20194 23418 20250 23420
rect 19954 23366 20000 23418
rect 20000 23366 20010 23418
rect 20034 23366 20064 23418
rect 20064 23366 20076 23418
rect 20076 23366 20090 23418
rect 20114 23366 20128 23418
rect 20128 23366 20140 23418
rect 20140 23366 20170 23418
rect 20194 23366 20204 23418
rect 20204 23366 20250 23418
rect 19954 23364 20010 23366
rect 20034 23364 20090 23366
rect 20114 23364 20170 23366
rect 20194 23364 20250 23366
rect 20626 25200 20682 25256
rect 19430 22652 19432 22672
rect 19432 22652 19484 22672
rect 19484 22652 19486 22672
rect 19430 22616 19486 22652
rect 20350 23024 20406 23080
rect 19338 21972 19340 21992
rect 19340 21972 19392 21992
rect 19392 21972 19394 21992
rect 19338 21936 19394 21972
rect 19430 21428 19432 21448
rect 19432 21428 19484 21448
rect 19484 21428 19486 21448
rect 19430 21392 19486 21428
rect 19706 22344 19762 22400
rect 19954 22330 20010 22332
rect 20034 22330 20090 22332
rect 20114 22330 20170 22332
rect 20194 22330 20250 22332
rect 19954 22278 20000 22330
rect 20000 22278 20010 22330
rect 20034 22278 20064 22330
rect 20064 22278 20076 22330
rect 20076 22278 20090 22330
rect 20114 22278 20128 22330
rect 20128 22278 20140 22330
rect 20140 22278 20170 22330
rect 20194 22278 20204 22330
rect 20204 22278 20250 22330
rect 19954 22276 20010 22278
rect 20034 22276 20090 22278
rect 20114 22276 20170 22278
rect 20194 22276 20250 22278
rect 19890 21972 19892 21992
rect 19892 21972 19944 21992
rect 19944 21972 19946 21992
rect 19890 21936 19946 21972
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 20534 22752 20590 22808
rect 20442 21936 20498 21992
rect 20902 22072 20958 22128
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 21638 26444 21694 26480
rect 21638 26424 21640 26444
rect 21640 26424 21692 26444
rect 21692 26424 21694 26444
rect 21454 24656 21510 24712
rect 21362 22888 21418 22944
rect 21362 20848 21418 20904
rect 21270 20576 21326 20632
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 6918 15544 6974 15600
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 21822 23704 21878 23760
rect 22668 27226 22724 27228
rect 22748 27226 22804 27228
rect 22828 27226 22884 27228
rect 22908 27226 22964 27228
rect 22668 27174 22714 27226
rect 22714 27174 22724 27226
rect 22748 27174 22778 27226
rect 22778 27174 22790 27226
rect 22790 27174 22804 27226
rect 22828 27174 22842 27226
rect 22842 27174 22854 27226
rect 22854 27174 22884 27226
rect 22908 27174 22918 27226
rect 22918 27174 22964 27226
rect 22668 27172 22724 27174
rect 22748 27172 22804 27174
rect 22828 27172 22884 27174
rect 22908 27172 22964 27174
rect 22668 26138 22724 26140
rect 22748 26138 22804 26140
rect 22828 26138 22884 26140
rect 22908 26138 22964 26140
rect 22668 26086 22714 26138
rect 22714 26086 22724 26138
rect 22748 26086 22778 26138
rect 22778 26086 22790 26138
rect 22790 26086 22804 26138
rect 22828 26086 22842 26138
rect 22842 26086 22854 26138
rect 22854 26086 22884 26138
rect 22908 26086 22918 26138
rect 22918 26086 22964 26138
rect 22668 26084 22724 26086
rect 22748 26084 22804 26086
rect 22828 26084 22884 26086
rect 22908 26084 22964 26086
rect 22668 25050 22724 25052
rect 22748 25050 22804 25052
rect 22828 25050 22884 25052
rect 22908 25050 22964 25052
rect 22668 24998 22714 25050
rect 22714 24998 22724 25050
rect 22748 24998 22778 25050
rect 22778 24998 22790 25050
rect 22790 24998 22804 25050
rect 22828 24998 22842 25050
rect 22842 24998 22854 25050
rect 22854 24998 22884 25050
rect 22908 24998 22918 25050
rect 22918 24998 22964 25050
rect 22668 24996 22724 24998
rect 22748 24996 22804 24998
rect 22828 24996 22884 24998
rect 22908 24996 22964 24998
rect 22668 23962 22724 23964
rect 22748 23962 22804 23964
rect 22828 23962 22884 23964
rect 22908 23962 22964 23964
rect 22668 23910 22714 23962
rect 22714 23910 22724 23962
rect 22748 23910 22778 23962
rect 22778 23910 22790 23962
rect 22790 23910 22804 23962
rect 22828 23910 22842 23962
rect 22842 23910 22854 23962
rect 22854 23910 22884 23962
rect 22908 23910 22918 23962
rect 22918 23910 22964 23962
rect 22668 23908 22724 23910
rect 22748 23908 22804 23910
rect 22828 23908 22884 23910
rect 22908 23908 22964 23910
rect 22190 23160 22246 23216
rect 22006 20304 22062 20360
rect 22006 19216 22062 19272
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 22006 16496 22062 16552
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 22668 22874 22724 22876
rect 22748 22874 22804 22876
rect 22828 22874 22884 22876
rect 22908 22874 22964 22876
rect 22668 22822 22714 22874
rect 22714 22822 22724 22874
rect 22748 22822 22778 22874
rect 22778 22822 22790 22874
rect 22790 22822 22804 22874
rect 22828 22822 22842 22874
rect 22842 22822 22854 22874
rect 22854 22822 22884 22874
rect 22908 22822 22918 22874
rect 22918 22822 22964 22874
rect 22668 22820 22724 22822
rect 22748 22820 22804 22822
rect 22828 22820 22884 22822
rect 22908 22820 22964 22822
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 22282 19760 22338 19816
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 22282 18708 22284 18728
rect 22284 18708 22336 18728
rect 22336 18708 22338 18728
rect 22282 18672 22338 18708
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 22282 18148 22338 18184
rect 22282 18128 22284 18148
rect 22284 18128 22336 18148
rect 22336 18128 22338 18148
rect 22282 17620 22284 17640
rect 22284 17620 22336 17640
rect 22336 17620 22338 17640
rect 22282 17584 22338 17620
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 22282 17060 22338 17096
rect 22282 17040 22284 17060
rect 22284 17040 22336 17060
rect 22336 17040 22338 17060
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 22098 15952 22154 16008
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 22282 15444 22284 15464
rect 22284 15444 22336 15464
rect 22336 15444 22338 15464
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 22282 15408 22338 15444
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 2870 11192 2926 11248
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 1582 10512 1638 10568
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 1582 9832 1638 9888
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 1582 9152 1638 9208
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 1766 8472 1822 8528
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 1582 7828 1584 7848
rect 1584 7828 1636 7848
rect 1636 7828 1638 7848
rect 1582 7792 1638 7828
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 22282 14884 22338 14920
rect 22282 14864 22284 14884
rect 22284 14864 22336 14884
rect 22336 14864 22338 14884
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 22282 13812 22284 13832
rect 22284 13812 22336 13832
rect 22336 13812 22338 13832
rect 22282 13776 22338 13812
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 22282 13268 22284 13288
rect 22284 13268 22336 13288
rect 22336 13268 22338 13288
rect 22282 13232 22338 13268
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 22282 12180 22284 12200
rect 22284 12180 22336 12200
rect 22336 12180 22338 12200
rect 22282 12144 22338 12180
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 22282 11620 22338 11656
rect 22282 11600 22284 11620
rect 22284 11600 22336 11620
rect 22336 11600 22338 11620
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 22282 10532 22338 10568
rect 22282 10512 22284 10532
rect 22284 10512 22336 10532
rect 22336 10512 22338 10532
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 22282 10004 22284 10024
rect 22284 10004 22336 10024
rect 22336 10004 22338 10024
rect 22282 9968 22338 10004
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 22282 8916 22284 8936
rect 22284 8916 22336 8936
rect 22336 8916 22338 8936
rect 22282 8880 22338 8916
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 22282 8356 22338 8392
rect 22282 8336 22284 8356
rect 22284 8336 22336 8356
rect 22336 8336 22338 8356
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 22282 7268 22338 7304
rect 22282 7248 22284 7268
rect 22284 7248 22336 7268
rect 22336 7248 22338 7268
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 22282 6740 22284 6760
rect 22284 6740 22336 6760
rect 22336 6740 22338 6760
rect 22282 6704 22338 6740
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 1674 5752 1730 5808
rect 22282 5652 22284 5672
rect 22284 5652 22336 5672
rect 22336 5652 22338 5672
rect 22282 5616 22338 5652
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 1582 5108 1584 5128
rect 1584 5108 1636 5128
rect 1636 5108 1638 5128
rect 1582 5072 1638 5108
rect 22282 5092 22338 5128
rect 22282 5072 22284 5092
rect 22284 5072 22336 5092
rect 22336 5072 22338 5092
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 22282 4004 22338 4040
rect 22282 3984 22284 4004
rect 22284 3984 22336 4004
rect 22336 3984 22338 4004
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 1582 3712 1638 3768
rect 22282 3476 22284 3496
rect 22284 3476 22336 3496
rect 22336 3476 22338 3496
rect 22282 3440 22338 3476
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 1582 3032 1638 3088
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
rect 1582 1672 1638 1728
rect 1398 992 1454 1048
<< metal3 >>
rect 0 28930 800 28960
rect 3969 28930 4035 28933
rect 0 28928 4035 28930
rect 0 28872 3974 28928
rect 4030 28872 4035 28928
rect 0 28870 4035 28872
rect 0 28840 800 28870
rect 3969 28867 4035 28870
rect 0 28250 800 28280
rect 4061 28250 4127 28253
rect 0 28248 4127 28250
rect 0 28192 4066 28248
rect 4122 28192 4127 28248
rect 0 28190 4127 28192
rect 0 28160 800 28190
rect 4061 28187 4127 28190
rect 3660 27776 3976 27777
rect 3660 27712 3666 27776
rect 3730 27712 3746 27776
rect 3810 27712 3826 27776
rect 3890 27712 3906 27776
rect 3970 27712 3976 27776
rect 3660 27711 3976 27712
rect 9088 27776 9404 27777
rect 9088 27712 9094 27776
rect 9158 27712 9174 27776
rect 9238 27712 9254 27776
rect 9318 27712 9334 27776
rect 9398 27712 9404 27776
rect 9088 27711 9404 27712
rect 14516 27776 14832 27777
rect 14516 27712 14522 27776
rect 14586 27712 14602 27776
rect 14666 27712 14682 27776
rect 14746 27712 14762 27776
rect 14826 27712 14832 27776
rect 14516 27711 14832 27712
rect 19944 27776 20260 27777
rect 19944 27712 19950 27776
rect 20014 27712 20030 27776
rect 20094 27712 20110 27776
rect 20174 27712 20190 27776
rect 20254 27712 20260 27776
rect 19944 27711 20260 27712
rect 0 27570 800 27600
rect 7189 27570 7255 27573
rect 0 27568 7255 27570
rect 0 27512 7194 27568
rect 7250 27512 7255 27568
rect 0 27510 7255 27512
rect 0 27480 800 27510
rect 7189 27507 7255 27510
rect 6374 27232 6690 27233
rect 6374 27168 6380 27232
rect 6444 27168 6460 27232
rect 6524 27168 6540 27232
rect 6604 27168 6620 27232
rect 6684 27168 6690 27232
rect 6374 27167 6690 27168
rect 11802 27232 12118 27233
rect 11802 27168 11808 27232
rect 11872 27168 11888 27232
rect 11952 27168 11968 27232
rect 12032 27168 12048 27232
rect 12112 27168 12118 27232
rect 11802 27167 12118 27168
rect 17230 27232 17546 27233
rect 17230 27168 17236 27232
rect 17300 27168 17316 27232
rect 17380 27168 17396 27232
rect 17460 27168 17476 27232
rect 17540 27168 17546 27232
rect 17230 27167 17546 27168
rect 22658 27232 22974 27233
rect 22658 27168 22664 27232
rect 22728 27168 22744 27232
rect 22808 27168 22824 27232
rect 22888 27168 22904 27232
rect 22968 27168 22974 27232
rect 22658 27167 22974 27168
rect 7005 27162 7071 27165
rect 8017 27162 8083 27165
rect 7005 27160 8083 27162
rect 7005 27104 7010 27160
rect 7066 27104 8022 27160
rect 8078 27104 8083 27160
rect 7005 27102 8083 27104
rect 7005 27099 7071 27102
rect 8017 27099 8083 27102
rect 5165 27026 5231 27029
rect 7281 27026 7347 27029
rect 7833 27026 7899 27029
rect 5165 27024 7899 27026
rect 5165 26968 5170 27024
rect 5226 26968 7286 27024
rect 7342 26968 7838 27024
rect 7894 26968 7899 27024
rect 5165 26966 7899 26968
rect 5165 26963 5231 26966
rect 7281 26963 7347 26966
rect 7833 26963 7899 26966
rect 0 26890 800 26920
rect 4061 26890 4127 26893
rect 0 26888 4127 26890
rect 0 26832 4066 26888
rect 4122 26832 4127 26888
rect 0 26830 4127 26832
rect 0 26800 800 26830
rect 4061 26827 4127 26830
rect 6729 26890 6795 26893
rect 7741 26890 7807 26893
rect 11237 26890 11303 26893
rect 6729 26888 11303 26890
rect 6729 26832 6734 26888
rect 6790 26832 7746 26888
rect 7802 26832 11242 26888
rect 11298 26832 11303 26888
rect 6729 26830 11303 26832
rect 6729 26827 6795 26830
rect 7741 26827 7807 26830
rect 11237 26827 11303 26830
rect 20529 26890 20595 26893
rect 23200 26890 24000 26920
rect 20529 26888 24000 26890
rect 20529 26832 20534 26888
rect 20590 26832 24000 26888
rect 20529 26830 24000 26832
rect 20529 26827 20595 26830
rect 23200 26800 24000 26830
rect 3660 26688 3976 26689
rect 3660 26624 3666 26688
rect 3730 26624 3746 26688
rect 3810 26624 3826 26688
rect 3890 26624 3906 26688
rect 3970 26624 3976 26688
rect 3660 26623 3976 26624
rect 9088 26688 9404 26689
rect 9088 26624 9094 26688
rect 9158 26624 9174 26688
rect 9238 26624 9254 26688
rect 9318 26624 9334 26688
rect 9398 26624 9404 26688
rect 9088 26623 9404 26624
rect 14516 26688 14832 26689
rect 14516 26624 14522 26688
rect 14586 26624 14602 26688
rect 14666 26624 14682 26688
rect 14746 26624 14762 26688
rect 14826 26624 14832 26688
rect 14516 26623 14832 26624
rect 19944 26688 20260 26689
rect 19944 26624 19950 26688
rect 20014 26624 20030 26688
rect 20094 26624 20110 26688
rect 20174 26624 20190 26688
rect 20254 26624 20260 26688
rect 19944 26623 20260 26624
rect 9765 26618 9831 26621
rect 11513 26618 11579 26621
rect 9765 26616 11579 26618
rect 9765 26560 9770 26616
rect 9826 26560 11518 26616
rect 11574 26560 11579 26616
rect 9765 26558 11579 26560
rect 9765 26555 9831 26558
rect 11513 26555 11579 26558
rect 6729 26482 6795 26485
rect 9857 26482 9923 26485
rect 6729 26480 9923 26482
rect 6729 26424 6734 26480
rect 6790 26424 9862 26480
rect 9918 26424 9923 26480
rect 6729 26422 9923 26424
rect 6729 26419 6795 26422
rect 9857 26419 9923 26422
rect 11973 26482 12039 26485
rect 14181 26482 14247 26485
rect 11973 26480 14247 26482
rect 11973 26424 11978 26480
rect 12034 26424 14186 26480
rect 14242 26424 14247 26480
rect 11973 26422 14247 26424
rect 11973 26419 12039 26422
rect 14181 26419 14247 26422
rect 21398 26420 21404 26484
rect 21468 26482 21474 26484
rect 21633 26482 21699 26485
rect 21468 26480 21699 26482
rect 21468 26424 21638 26480
rect 21694 26424 21699 26480
rect 21468 26422 21699 26424
rect 21468 26420 21474 26422
rect 21633 26419 21699 26422
rect 2957 26346 3023 26349
rect 4102 26346 4108 26348
rect 2957 26344 4108 26346
rect 2957 26288 2962 26344
rect 3018 26288 4108 26344
rect 2957 26286 4108 26288
rect 2957 26283 3023 26286
rect 4102 26284 4108 26286
rect 4172 26284 4178 26348
rect 5349 26346 5415 26349
rect 8293 26346 8359 26349
rect 5349 26344 8359 26346
rect 5349 26288 5354 26344
rect 5410 26288 8298 26344
rect 8354 26288 8359 26344
rect 5349 26286 8359 26288
rect 5349 26283 5415 26286
rect 8293 26283 8359 26286
rect 9121 26346 9187 26349
rect 11329 26346 11395 26349
rect 14273 26346 14339 26349
rect 9121 26344 14339 26346
rect 9121 26288 9126 26344
rect 9182 26288 11334 26344
rect 11390 26288 14278 26344
rect 14334 26288 14339 26344
rect 9121 26286 14339 26288
rect 9121 26283 9187 26286
rect 11329 26283 11395 26286
rect 14273 26283 14339 26286
rect 19425 26346 19491 26349
rect 23200 26346 24000 26376
rect 19425 26344 24000 26346
rect 19425 26288 19430 26344
rect 19486 26288 24000 26344
rect 19425 26286 24000 26288
rect 19425 26283 19491 26286
rect 23200 26256 24000 26286
rect 0 26210 800 26240
rect 4061 26210 4127 26213
rect 0 26208 4127 26210
rect 0 26152 4066 26208
rect 4122 26152 4127 26208
rect 0 26150 4127 26152
rect 0 26120 800 26150
rect 4061 26147 4127 26150
rect 6374 26144 6690 26145
rect 6374 26080 6380 26144
rect 6444 26080 6460 26144
rect 6524 26080 6540 26144
rect 6604 26080 6620 26144
rect 6684 26080 6690 26144
rect 6374 26079 6690 26080
rect 11802 26144 12118 26145
rect 11802 26080 11808 26144
rect 11872 26080 11888 26144
rect 11952 26080 11968 26144
rect 12032 26080 12048 26144
rect 12112 26080 12118 26144
rect 11802 26079 12118 26080
rect 17230 26144 17546 26145
rect 17230 26080 17236 26144
rect 17300 26080 17316 26144
rect 17380 26080 17396 26144
rect 17460 26080 17476 26144
rect 17540 26080 17546 26144
rect 17230 26079 17546 26080
rect 22658 26144 22974 26145
rect 22658 26080 22664 26144
rect 22728 26080 22744 26144
rect 22808 26080 22824 26144
rect 22888 26080 22904 26144
rect 22968 26080 22974 26144
rect 22658 26079 22974 26080
rect 9673 25938 9739 25941
rect 10501 25938 10567 25941
rect 9673 25936 10567 25938
rect 9673 25880 9678 25936
rect 9734 25880 10506 25936
rect 10562 25880 10567 25936
rect 9673 25878 10567 25880
rect 9673 25875 9739 25878
rect 10501 25875 10567 25878
rect 7833 25802 7899 25805
rect 12893 25802 12959 25805
rect 7833 25800 12959 25802
rect 7833 25744 7838 25800
rect 7894 25744 12898 25800
rect 12954 25744 12959 25800
rect 7833 25742 12959 25744
rect 7833 25739 7899 25742
rect 12893 25739 12959 25742
rect 13077 25802 13143 25805
rect 14365 25802 14431 25805
rect 13077 25800 14431 25802
rect 13077 25744 13082 25800
rect 13138 25744 14370 25800
rect 14426 25744 14431 25800
rect 13077 25742 14431 25744
rect 13077 25739 13143 25742
rect 14365 25739 14431 25742
rect 19425 25802 19491 25805
rect 23200 25802 24000 25832
rect 19425 25800 24000 25802
rect 19425 25744 19430 25800
rect 19486 25744 24000 25800
rect 19425 25742 24000 25744
rect 19425 25739 19491 25742
rect 23200 25712 24000 25742
rect 3660 25600 3976 25601
rect 0 25530 800 25560
rect 3660 25536 3666 25600
rect 3730 25536 3746 25600
rect 3810 25536 3826 25600
rect 3890 25536 3906 25600
rect 3970 25536 3976 25600
rect 3660 25535 3976 25536
rect 9088 25600 9404 25601
rect 9088 25536 9094 25600
rect 9158 25536 9174 25600
rect 9238 25536 9254 25600
rect 9318 25536 9334 25600
rect 9398 25536 9404 25600
rect 9088 25535 9404 25536
rect 14516 25600 14832 25601
rect 14516 25536 14522 25600
rect 14586 25536 14602 25600
rect 14666 25536 14682 25600
rect 14746 25536 14762 25600
rect 14826 25536 14832 25600
rect 14516 25535 14832 25536
rect 19944 25600 20260 25601
rect 19944 25536 19950 25600
rect 20014 25536 20030 25600
rect 20094 25536 20110 25600
rect 20174 25536 20190 25600
rect 20254 25536 20260 25600
rect 19944 25535 20260 25536
rect 3417 25530 3483 25533
rect 0 25528 3483 25530
rect 0 25472 3422 25528
rect 3478 25472 3483 25528
rect 0 25470 3483 25472
rect 0 25440 800 25470
rect 3417 25467 3483 25470
rect 1209 25394 1275 25397
rect 6269 25394 6335 25397
rect 1209 25392 6335 25394
rect 1209 25336 1214 25392
rect 1270 25336 6274 25392
rect 6330 25336 6335 25392
rect 1209 25334 6335 25336
rect 1209 25331 1275 25334
rect 6269 25331 6335 25334
rect 20621 25258 20687 25261
rect 23200 25258 24000 25288
rect 20621 25256 24000 25258
rect 20621 25200 20626 25256
rect 20682 25200 24000 25256
rect 20621 25198 24000 25200
rect 20621 25195 20687 25198
rect 23200 25168 24000 25198
rect 6374 25056 6690 25057
rect 6374 24992 6380 25056
rect 6444 24992 6460 25056
rect 6524 24992 6540 25056
rect 6604 24992 6620 25056
rect 6684 24992 6690 25056
rect 6374 24991 6690 24992
rect 11802 25056 12118 25057
rect 11802 24992 11808 25056
rect 11872 24992 11888 25056
rect 11952 24992 11968 25056
rect 12032 24992 12048 25056
rect 12112 24992 12118 25056
rect 11802 24991 12118 24992
rect 17230 25056 17546 25057
rect 17230 24992 17236 25056
rect 17300 24992 17316 25056
rect 17380 24992 17396 25056
rect 17460 24992 17476 25056
rect 17540 24992 17546 25056
rect 17230 24991 17546 24992
rect 22658 25056 22974 25057
rect 22658 24992 22664 25056
rect 22728 24992 22744 25056
rect 22808 24992 22824 25056
rect 22888 24992 22904 25056
rect 22968 24992 22974 25056
rect 22658 24991 22974 24992
rect 4286 24924 4292 24988
rect 4356 24986 4362 24988
rect 5073 24986 5139 24989
rect 4356 24984 5139 24986
rect 4356 24928 5078 24984
rect 5134 24928 5139 24984
rect 4356 24926 5139 24928
rect 4356 24924 4362 24926
rect 5073 24923 5139 24926
rect 0 24850 800 24880
rect 2497 24850 2563 24853
rect 0 24848 2563 24850
rect 0 24792 2502 24848
rect 2558 24792 2563 24848
rect 0 24790 2563 24792
rect 0 24760 800 24790
rect 2497 24787 2563 24790
rect 2681 24714 2747 24717
rect 5349 24714 5415 24717
rect 2681 24712 5415 24714
rect 2681 24656 2686 24712
rect 2742 24656 5354 24712
rect 5410 24656 5415 24712
rect 2681 24654 5415 24656
rect 2681 24651 2747 24654
rect 5349 24651 5415 24654
rect 21449 24714 21515 24717
rect 23200 24714 24000 24744
rect 21449 24712 24000 24714
rect 21449 24656 21454 24712
rect 21510 24656 24000 24712
rect 21449 24654 24000 24656
rect 21449 24651 21515 24654
rect 23200 24624 24000 24654
rect 3660 24512 3976 24513
rect 3660 24448 3666 24512
rect 3730 24448 3746 24512
rect 3810 24448 3826 24512
rect 3890 24448 3906 24512
rect 3970 24448 3976 24512
rect 3660 24447 3976 24448
rect 9088 24512 9404 24513
rect 9088 24448 9094 24512
rect 9158 24448 9174 24512
rect 9238 24448 9254 24512
rect 9318 24448 9334 24512
rect 9398 24448 9404 24512
rect 9088 24447 9404 24448
rect 14516 24512 14832 24513
rect 14516 24448 14522 24512
rect 14586 24448 14602 24512
rect 14666 24448 14682 24512
rect 14746 24448 14762 24512
rect 14826 24448 14832 24512
rect 14516 24447 14832 24448
rect 19944 24512 20260 24513
rect 19944 24448 19950 24512
rect 20014 24448 20030 24512
rect 20094 24448 20110 24512
rect 20174 24448 20190 24512
rect 20254 24448 20260 24512
rect 19944 24447 20260 24448
rect 2681 24306 2747 24309
rect 6637 24306 6703 24309
rect 2681 24304 6703 24306
rect 2681 24248 2686 24304
rect 2742 24248 6642 24304
rect 6698 24248 6703 24304
rect 2681 24246 6703 24248
rect 2681 24243 2747 24246
rect 6637 24243 6703 24246
rect 0 24170 800 24200
rect 4061 24170 4127 24173
rect 0 24168 4127 24170
rect 0 24112 4066 24168
rect 4122 24112 4127 24168
rect 0 24110 4127 24112
rect 0 24080 800 24110
rect 4061 24107 4127 24110
rect 19333 24170 19399 24173
rect 23200 24170 24000 24200
rect 19333 24168 24000 24170
rect 19333 24112 19338 24168
rect 19394 24112 24000 24168
rect 19333 24110 24000 24112
rect 19333 24107 19399 24110
rect 23200 24080 24000 24110
rect 2589 24034 2655 24037
rect 5165 24034 5231 24037
rect 2589 24032 5231 24034
rect 2589 23976 2594 24032
rect 2650 23976 5170 24032
rect 5226 23976 5231 24032
rect 2589 23974 5231 23976
rect 2589 23971 2655 23974
rect 5165 23971 5231 23974
rect 5168 23762 5228 23971
rect 6374 23968 6690 23969
rect 6374 23904 6380 23968
rect 6444 23904 6460 23968
rect 6524 23904 6540 23968
rect 6604 23904 6620 23968
rect 6684 23904 6690 23968
rect 6374 23903 6690 23904
rect 11802 23968 12118 23969
rect 11802 23904 11808 23968
rect 11872 23904 11888 23968
rect 11952 23904 11968 23968
rect 12032 23904 12048 23968
rect 12112 23904 12118 23968
rect 11802 23903 12118 23904
rect 17230 23968 17546 23969
rect 17230 23904 17236 23968
rect 17300 23904 17316 23968
rect 17380 23904 17396 23968
rect 17460 23904 17476 23968
rect 17540 23904 17546 23968
rect 17230 23903 17546 23904
rect 22658 23968 22974 23969
rect 22658 23904 22664 23968
rect 22728 23904 22744 23968
rect 22808 23904 22824 23968
rect 22888 23904 22904 23968
rect 22968 23904 22974 23968
rect 22658 23903 22974 23904
rect 6729 23762 6795 23765
rect 5168 23760 6795 23762
rect 5168 23704 6734 23760
rect 6790 23704 6795 23760
rect 5168 23702 6795 23704
rect 6729 23699 6795 23702
rect 19425 23762 19491 23765
rect 21817 23762 21883 23765
rect 19425 23760 21883 23762
rect 19425 23704 19430 23760
rect 19486 23704 21822 23760
rect 21878 23704 21883 23760
rect 19425 23702 21883 23704
rect 19425 23699 19491 23702
rect 21817 23699 21883 23702
rect 3601 23626 3667 23629
rect 5257 23626 5323 23629
rect 3601 23624 5323 23626
rect 3601 23568 3606 23624
rect 3662 23568 5262 23624
rect 5318 23568 5323 23624
rect 3601 23566 5323 23568
rect 3601 23563 3667 23566
rect 5257 23563 5323 23566
rect 19793 23626 19859 23629
rect 23200 23626 24000 23656
rect 19793 23624 24000 23626
rect 19793 23568 19798 23624
rect 19854 23568 24000 23624
rect 19793 23566 24000 23568
rect 19793 23563 19859 23566
rect 23200 23536 24000 23566
rect 0 23490 800 23520
rect 2865 23490 2931 23493
rect 0 23488 2931 23490
rect 0 23432 2870 23488
rect 2926 23432 2931 23488
rect 0 23430 2931 23432
rect 0 23400 800 23430
rect 2865 23427 2931 23430
rect 3660 23424 3976 23425
rect 3660 23360 3666 23424
rect 3730 23360 3746 23424
rect 3810 23360 3826 23424
rect 3890 23360 3906 23424
rect 3970 23360 3976 23424
rect 3660 23359 3976 23360
rect 9088 23424 9404 23425
rect 9088 23360 9094 23424
rect 9158 23360 9174 23424
rect 9238 23360 9254 23424
rect 9318 23360 9334 23424
rect 9398 23360 9404 23424
rect 9088 23359 9404 23360
rect 14516 23424 14832 23425
rect 14516 23360 14522 23424
rect 14586 23360 14602 23424
rect 14666 23360 14682 23424
rect 14746 23360 14762 23424
rect 14826 23360 14832 23424
rect 14516 23359 14832 23360
rect 19944 23424 20260 23425
rect 19944 23360 19950 23424
rect 20014 23360 20030 23424
rect 20094 23360 20110 23424
rect 20174 23360 20190 23424
rect 20254 23360 20260 23424
rect 19944 23359 20260 23360
rect 4153 23220 4219 23221
rect 4102 23218 4108 23220
rect 4062 23158 4108 23218
rect 4172 23216 4219 23220
rect 4214 23160 4219 23216
rect 4102 23156 4108 23158
rect 4172 23156 4219 23160
rect 4153 23155 4219 23156
rect 4337 23218 4403 23221
rect 4797 23218 4863 23221
rect 4337 23216 4863 23218
rect 4337 23160 4342 23216
rect 4398 23160 4802 23216
rect 4858 23160 4863 23216
rect 4337 23158 4863 23160
rect 4337 23155 4403 23158
rect 4797 23155 4863 23158
rect 17033 23218 17099 23221
rect 22185 23218 22251 23221
rect 17033 23216 22251 23218
rect 17033 23160 17038 23216
rect 17094 23160 22190 23216
rect 22246 23160 22251 23216
rect 17033 23158 22251 23160
rect 17033 23155 17099 23158
rect 22185 23155 22251 23158
rect 20345 23082 20411 23085
rect 23200 23082 24000 23112
rect 20345 23080 24000 23082
rect 20345 23024 20350 23080
rect 20406 23024 24000 23080
rect 20345 23022 24000 23024
rect 20345 23019 20411 23022
rect 23200 22992 24000 23022
rect 19517 22946 19583 22949
rect 21357 22946 21423 22949
rect 19517 22944 21423 22946
rect 19517 22888 19522 22944
rect 19578 22888 21362 22944
rect 21418 22888 21423 22944
rect 19517 22886 21423 22888
rect 19517 22883 19583 22886
rect 21357 22883 21423 22886
rect 6374 22880 6690 22881
rect 0 22810 800 22840
rect 6374 22816 6380 22880
rect 6444 22816 6460 22880
rect 6524 22816 6540 22880
rect 6604 22816 6620 22880
rect 6684 22816 6690 22880
rect 6374 22815 6690 22816
rect 11802 22880 12118 22881
rect 11802 22816 11808 22880
rect 11872 22816 11888 22880
rect 11952 22816 11968 22880
rect 12032 22816 12048 22880
rect 12112 22816 12118 22880
rect 11802 22815 12118 22816
rect 17230 22880 17546 22881
rect 17230 22816 17236 22880
rect 17300 22816 17316 22880
rect 17380 22816 17396 22880
rect 17460 22816 17476 22880
rect 17540 22816 17546 22880
rect 17230 22815 17546 22816
rect 22658 22880 22974 22881
rect 22658 22816 22664 22880
rect 22728 22816 22744 22880
rect 22808 22816 22824 22880
rect 22888 22816 22904 22880
rect 22968 22816 22974 22880
rect 22658 22815 22974 22816
rect 4061 22810 4127 22813
rect 20529 22810 20595 22813
rect 0 22808 4127 22810
rect 0 22752 4066 22808
rect 4122 22752 4127 22808
rect 0 22750 4127 22752
rect 0 22720 800 22750
rect 4061 22747 4127 22750
rect 19428 22808 20595 22810
rect 19428 22752 20534 22808
rect 20590 22752 20595 22808
rect 19428 22750 20595 22752
rect 19428 22677 19488 22750
rect 20529 22747 20595 22750
rect 19425 22672 19491 22677
rect 19425 22616 19430 22672
rect 19486 22616 19491 22672
rect 19425 22611 19491 22616
rect 3877 22538 3943 22541
rect 23200 22538 24000 22568
rect 2730 22536 3943 22538
rect 2730 22480 3882 22536
rect 3938 22480 3943 22536
rect 2730 22478 3943 22480
rect 0 22130 800 22160
rect 2730 22130 2790 22478
rect 3877 22475 3943 22478
rect 19750 22478 24000 22538
rect 19750 22405 19810 22478
rect 23200 22448 24000 22478
rect 19701 22400 19810 22405
rect 19701 22344 19706 22400
rect 19762 22344 19810 22400
rect 19701 22342 19810 22344
rect 19701 22339 19767 22342
rect 3660 22336 3976 22337
rect 3660 22272 3666 22336
rect 3730 22272 3746 22336
rect 3810 22272 3826 22336
rect 3890 22272 3906 22336
rect 3970 22272 3976 22336
rect 3660 22271 3976 22272
rect 9088 22336 9404 22337
rect 9088 22272 9094 22336
rect 9158 22272 9174 22336
rect 9238 22272 9254 22336
rect 9318 22272 9334 22336
rect 9398 22272 9404 22336
rect 9088 22271 9404 22272
rect 14516 22336 14832 22337
rect 14516 22272 14522 22336
rect 14586 22272 14602 22336
rect 14666 22272 14682 22336
rect 14746 22272 14762 22336
rect 14826 22272 14832 22336
rect 14516 22271 14832 22272
rect 19944 22336 20260 22337
rect 19944 22272 19950 22336
rect 20014 22272 20030 22336
rect 20094 22272 20110 22336
rect 20174 22272 20190 22336
rect 20254 22272 20260 22336
rect 19944 22271 20260 22272
rect 0 22070 2790 22130
rect 3877 22130 3943 22133
rect 5441 22130 5507 22133
rect 3877 22128 5507 22130
rect 3877 22072 3882 22128
rect 3938 22072 5446 22128
rect 5502 22072 5507 22128
rect 3877 22070 5507 22072
rect 0 22040 800 22070
rect 3877 22067 3943 22070
rect 5441 22067 5507 22070
rect 17585 22130 17651 22133
rect 20897 22130 20963 22133
rect 17585 22128 20963 22130
rect 17585 22072 17590 22128
rect 17646 22072 20902 22128
rect 20958 22072 20963 22128
rect 17585 22070 20963 22072
rect 17585 22067 17651 22070
rect 20897 22067 20963 22070
rect 19333 21994 19399 21997
rect 19885 21994 19951 21997
rect 19333 21992 19951 21994
rect 19333 21936 19338 21992
rect 19394 21936 19890 21992
rect 19946 21936 19951 21992
rect 19333 21934 19951 21936
rect 19333 21931 19399 21934
rect 19885 21931 19951 21934
rect 20437 21994 20503 21997
rect 23200 21994 24000 22024
rect 20437 21992 24000 21994
rect 20437 21936 20442 21992
rect 20498 21936 24000 21992
rect 20437 21934 24000 21936
rect 20437 21931 20503 21934
rect 23200 21904 24000 21934
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 2129 21722 2195 21725
rect 4286 21722 4292 21724
rect 2129 21720 4292 21722
rect 2129 21664 2134 21720
rect 2190 21664 4292 21720
rect 2129 21662 4292 21664
rect 2129 21659 2195 21662
rect 4286 21660 4292 21662
rect 4356 21660 4362 21724
rect 0 21450 800 21480
rect 3141 21450 3207 21453
rect 0 21448 3207 21450
rect 0 21392 3146 21448
rect 3202 21392 3207 21448
rect 0 21390 3207 21392
rect 0 21360 800 21390
rect 3141 21387 3207 21390
rect 19425 21450 19491 21453
rect 23200 21450 24000 21480
rect 19425 21448 24000 21450
rect 19425 21392 19430 21448
rect 19486 21392 24000 21448
rect 19425 21390 24000 21392
rect 19425 21387 19491 21390
rect 23200 21360 24000 21390
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 21357 20906 21423 20909
rect 23200 20906 24000 20936
rect 21357 20904 24000 20906
rect 21357 20848 21362 20904
rect 21418 20848 24000 20904
rect 21357 20846 24000 20848
rect 21357 20843 21423 20846
rect 23200 20816 24000 20846
rect 0 20770 800 20800
rect 3049 20770 3115 20773
rect 0 20768 3115 20770
rect 0 20712 3054 20768
rect 3110 20712 3115 20768
rect 0 20710 3115 20712
rect 0 20680 800 20710
rect 3049 20707 3115 20710
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 21265 20634 21331 20637
rect 21398 20634 21404 20636
rect 21265 20632 21404 20634
rect 21265 20576 21270 20632
rect 21326 20576 21404 20632
rect 21265 20574 21404 20576
rect 21265 20571 21331 20574
rect 21398 20572 21404 20574
rect 21468 20572 21474 20636
rect 22001 20362 22067 20365
rect 23200 20362 24000 20392
rect 22001 20360 24000 20362
rect 22001 20304 22006 20360
rect 22062 20304 24000 20360
rect 22001 20302 24000 20304
rect 22001 20299 22067 20302
rect 23200 20272 24000 20302
rect 3660 20160 3976 20161
rect 0 20090 800 20120
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 2405 20090 2471 20093
rect 0 20088 2471 20090
rect 0 20032 2410 20088
rect 2466 20032 2471 20088
rect 0 20030 2471 20032
rect 0 20000 800 20030
rect 2405 20027 2471 20030
rect 22277 19818 22343 19821
rect 23200 19818 24000 19848
rect 22277 19816 24000 19818
rect 22277 19760 22282 19816
rect 22338 19760 24000 19816
rect 22277 19758 24000 19760
rect 22277 19755 22343 19758
rect 23200 19728 24000 19758
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 0 19410 800 19440
rect 2221 19410 2287 19413
rect 0 19408 2287 19410
rect 0 19352 2226 19408
rect 2282 19352 2287 19408
rect 0 19350 2287 19352
rect 0 19320 800 19350
rect 2221 19347 2287 19350
rect 2405 19410 2471 19413
rect 5022 19410 5028 19412
rect 2405 19408 5028 19410
rect 2405 19352 2410 19408
rect 2466 19352 5028 19408
rect 2405 19350 5028 19352
rect 2405 19347 2471 19350
rect 5022 19348 5028 19350
rect 5092 19348 5098 19412
rect 22001 19274 22067 19277
rect 23200 19274 24000 19304
rect 22001 19272 24000 19274
rect 22001 19216 22006 19272
rect 22062 19216 24000 19272
rect 22001 19214 24000 19216
rect 22001 19211 22067 19214
rect 23200 19184 24000 19214
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 22277 18730 22343 18733
rect 23200 18730 24000 18760
rect 22277 18728 24000 18730
rect 22277 18672 22282 18728
rect 22338 18672 24000 18728
rect 22277 18670 24000 18672
rect 22277 18667 22343 18670
rect 23200 18640 24000 18670
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 1945 18186 2011 18189
rect 4286 18186 4292 18188
rect 1945 18184 4292 18186
rect 1945 18128 1950 18184
rect 2006 18128 4292 18184
rect 1945 18126 4292 18128
rect 1945 18123 2011 18126
rect 4286 18124 4292 18126
rect 4356 18124 4362 18188
rect 22277 18186 22343 18189
rect 23200 18186 24000 18216
rect 22277 18184 24000 18186
rect 22277 18128 22282 18184
rect 22338 18128 24000 18184
rect 22277 18126 24000 18128
rect 22277 18123 22343 18126
rect 23200 18096 24000 18126
rect 0 18050 800 18080
rect 3509 18050 3575 18053
rect 0 18048 3575 18050
rect 0 17992 3514 18048
rect 3570 17992 3575 18048
rect 0 17990 3575 17992
rect 0 17960 800 17990
rect 3509 17987 3575 17990
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 22277 17642 22343 17645
rect 23200 17642 24000 17672
rect 22277 17640 24000 17642
rect 22277 17584 22282 17640
rect 22338 17584 24000 17640
rect 22277 17582 24000 17584
rect 22277 17579 22343 17582
rect 23200 17552 24000 17582
rect 6374 17440 6690 17441
rect 0 17370 800 17400
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 22277 17098 22343 17101
rect 23200 17098 24000 17128
rect 22277 17096 24000 17098
rect 22277 17040 22282 17096
rect 22338 17040 24000 17096
rect 22277 17038 24000 17040
rect 22277 17035 22343 17038
rect 23200 17008 24000 17038
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 0 16690 800 16720
rect 2773 16690 2839 16693
rect 0 16688 2839 16690
rect 0 16632 2778 16688
rect 2834 16632 2839 16688
rect 0 16630 2839 16632
rect 0 16600 800 16630
rect 2773 16627 2839 16630
rect 22001 16554 22067 16557
rect 23200 16554 24000 16584
rect 22001 16552 24000 16554
rect 22001 16496 22006 16552
rect 22062 16496 24000 16552
rect 22001 16494 24000 16496
rect 22001 16491 22067 16494
rect 23200 16464 24000 16494
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 0 16010 800 16040
rect 4153 16010 4219 16013
rect 0 16008 4219 16010
rect 0 15952 4158 16008
rect 4214 15952 4219 16008
rect 0 15950 4219 15952
rect 0 15920 800 15950
rect 4153 15947 4219 15950
rect 22093 16010 22159 16013
rect 23200 16010 24000 16040
rect 22093 16008 24000 16010
rect 22093 15952 22098 16008
rect 22154 15952 24000 16008
rect 22093 15950 24000 15952
rect 22093 15947 22159 15950
rect 23200 15920 24000 15950
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 5073 15740 5139 15741
rect 5022 15676 5028 15740
rect 5092 15738 5139 15740
rect 5092 15736 5184 15738
rect 5134 15680 5184 15736
rect 5092 15678 5184 15680
rect 5092 15676 5139 15678
rect 5073 15675 5139 15676
rect 2681 15602 2747 15605
rect 3049 15602 3115 15605
rect 4337 15602 4403 15605
rect 6913 15602 6979 15605
rect 2681 15600 6979 15602
rect 2681 15544 2686 15600
rect 2742 15544 3054 15600
rect 3110 15544 4342 15600
rect 4398 15544 6918 15600
rect 6974 15544 6979 15600
rect 2681 15542 6979 15544
rect 2681 15539 2747 15542
rect 3049 15539 3115 15542
rect 4337 15539 4403 15542
rect 6913 15539 6979 15542
rect 22277 15466 22343 15469
rect 23200 15466 24000 15496
rect 22277 15464 24000 15466
rect 22277 15408 22282 15464
rect 22338 15408 24000 15464
rect 22277 15406 24000 15408
rect 22277 15403 22343 15406
rect 23200 15376 24000 15406
rect 0 15330 800 15360
rect 3049 15330 3115 15333
rect 0 15328 3115 15330
rect 0 15272 3054 15328
rect 3110 15272 3115 15328
rect 0 15270 3115 15272
rect 0 15240 800 15270
rect 3049 15267 3115 15270
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 3601 14922 3667 14925
rect 3374 14920 3667 14922
rect 3374 14864 3606 14920
rect 3662 14864 3667 14920
rect 3374 14862 3667 14864
rect 3374 14789 3434 14862
rect 3601 14859 3667 14862
rect 22277 14922 22343 14925
rect 23200 14922 24000 14952
rect 22277 14920 24000 14922
rect 22277 14864 22282 14920
rect 22338 14864 24000 14920
rect 22277 14862 24000 14864
rect 22277 14859 22343 14862
rect 23200 14832 24000 14862
rect 3325 14784 3434 14789
rect 3325 14728 3330 14784
rect 3386 14728 3434 14784
rect 3325 14726 3434 14728
rect 3325 14723 3391 14726
rect 3660 14720 3976 14721
rect 0 14650 800 14680
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 0 14590 2790 14650
rect 0 14560 800 14590
rect 2730 14378 2790 14590
rect 4337 14516 4403 14517
rect 4286 14452 4292 14516
rect 4356 14514 4403 14516
rect 4356 14512 4448 14514
rect 4398 14456 4448 14512
rect 4356 14454 4448 14456
rect 4356 14452 4403 14454
rect 4337 14451 4403 14452
rect 3509 14378 3575 14381
rect 2730 14376 3575 14378
rect 2730 14320 3514 14376
rect 3570 14320 3575 14376
rect 2730 14318 3575 14320
rect 3509 14315 3575 14318
rect 23200 14288 24000 14408
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 0 13970 800 14000
rect 3877 13970 3943 13973
rect 0 13968 3943 13970
rect 0 13912 3882 13968
rect 3938 13912 3943 13968
rect 0 13910 3943 13912
rect 0 13880 800 13910
rect 3877 13907 3943 13910
rect 22277 13834 22343 13837
rect 23200 13834 24000 13864
rect 22277 13832 24000 13834
rect 22277 13776 22282 13832
rect 22338 13776 24000 13832
rect 22277 13774 24000 13776
rect 22277 13771 22343 13774
rect 23200 13744 24000 13774
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 0 13290 800 13320
rect 2773 13290 2839 13293
rect 0 13288 2839 13290
rect 0 13232 2778 13288
rect 2834 13232 2839 13288
rect 0 13230 2839 13232
rect 0 13200 800 13230
rect 2773 13227 2839 13230
rect 22277 13290 22343 13293
rect 23200 13290 24000 13320
rect 22277 13288 24000 13290
rect 22277 13232 22282 13288
rect 22338 13232 24000 13288
rect 22277 13230 24000 13232
rect 22277 13227 22343 13230
rect 23200 13200 24000 13230
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 23200 12656 24000 12776
rect 0 12610 800 12640
rect 3509 12610 3575 12613
rect 0 12608 3575 12610
rect 0 12552 3514 12608
rect 3570 12552 3575 12608
rect 0 12550 3575 12552
rect 0 12520 800 12550
rect 3509 12547 3575 12550
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 22277 12202 22343 12205
rect 23200 12202 24000 12232
rect 22277 12200 24000 12202
rect 22277 12144 22282 12200
rect 22338 12144 24000 12200
rect 22277 12142 24000 12144
rect 22277 12139 22343 12142
rect 23200 12112 24000 12142
rect 6374 12000 6690 12001
rect 0 11930 800 11960
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 2221 11930 2287 11933
rect 0 11928 2287 11930
rect 0 11872 2226 11928
rect 2282 11872 2287 11928
rect 0 11870 2287 11872
rect 0 11840 800 11870
rect 2221 11867 2287 11870
rect 22277 11658 22343 11661
rect 23200 11658 24000 11688
rect 22277 11656 24000 11658
rect 22277 11600 22282 11656
rect 22338 11600 24000 11656
rect 22277 11598 24000 11600
rect 22277 11595 22343 11598
rect 23200 11568 24000 11598
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 0 11250 800 11280
rect 2865 11250 2931 11253
rect 0 11248 2931 11250
rect 0 11192 2870 11248
rect 2926 11192 2931 11248
rect 0 11190 2931 11192
rect 0 11160 800 11190
rect 2865 11187 2931 11190
rect 23200 11024 24000 11144
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 0 10570 800 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 800 10510
rect 1577 10507 1643 10510
rect 22277 10570 22343 10573
rect 23200 10570 24000 10600
rect 22277 10568 24000 10570
rect 22277 10512 22282 10568
rect 22338 10512 24000 10568
rect 22277 10510 24000 10512
rect 22277 10507 22343 10510
rect 23200 10480 24000 10510
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 22277 10026 22343 10029
rect 23200 10026 24000 10056
rect 22277 10024 24000 10026
rect 22277 9968 22282 10024
rect 22338 9968 24000 10024
rect 22277 9966 24000 9968
rect 22277 9963 22343 9966
rect 23200 9936 24000 9966
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 23200 9392 24000 9512
rect 3660 9280 3976 9281
rect 0 9210 800 9240
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 22277 8938 22343 8941
rect 23200 8938 24000 8968
rect 22277 8936 24000 8938
rect 22277 8880 22282 8936
rect 22338 8880 24000 8936
rect 22277 8878 24000 8880
rect 22277 8875 22343 8878
rect 23200 8848 24000 8878
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 0 8530 800 8560
rect 1761 8530 1827 8533
rect 0 8528 1827 8530
rect 0 8472 1766 8528
rect 1822 8472 1827 8528
rect 0 8470 1827 8472
rect 0 8440 800 8470
rect 1761 8467 1827 8470
rect 22277 8394 22343 8397
rect 23200 8394 24000 8424
rect 22277 8392 24000 8394
rect 22277 8336 22282 8392
rect 22338 8336 24000 8392
rect 22277 8334 24000 8336
rect 22277 8331 22343 8334
rect 23200 8304 24000 8334
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 23200 7760 24000 7880
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 22277 7306 22343 7309
rect 23200 7306 24000 7336
rect 22277 7304 24000 7306
rect 22277 7248 22282 7304
rect 22338 7248 24000 7304
rect 22277 7246 24000 7248
rect 22277 7243 22343 7246
rect 23200 7216 24000 7246
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 22277 6762 22343 6765
rect 23200 6762 24000 6792
rect 22277 6760 24000 6762
rect 22277 6704 22282 6760
rect 22338 6704 24000 6760
rect 22277 6702 24000 6704
rect 22277 6699 22343 6702
rect 23200 6672 24000 6702
rect 6374 6560 6690 6561
rect 0 6400 800 6520
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 23200 6128 24000 6248
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 22277 5674 22343 5677
rect 23200 5674 24000 5704
rect 22277 5672 24000 5674
rect 22277 5616 22282 5672
rect 22338 5616 24000 5672
rect 22277 5614 24000 5616
rect 22277 5611 22343 5614
rect 23200 5584 24000 5614
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 22277 5130 22343 5133
rect 23200 5130 24000 5160
rect 22277 5128 24000 5130
rect 22277 5072 22282 5128
rect 22338 5072 24000 5128
rect 22277 5070 24000 5072
rect 22277 5067 22343 5070
rect 23200 5040 24000 5070
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 23200 4496 24000 4616
rect 0 4360 800 4480
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 22277 4042 22343 4045
rect 23200 4042 24000 4072
rect 22277 4040 24000 4042
rect 22277 3984 22282 4040
rect 22338 3984 24000 4040
rect 22277 3982 24000 3984
rect 22277 3979 22343 3982
rect 23200 3952 24000 3982
rect 3660 3840 3976 3841
rect 0 3770 800 3800
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 22277 3498 22343 3501
rect 23200 3498 24000 3528
rect 22277 3496 24000 3498
rect 22277 3440 22282 3496
rect 22338 3440 24000 3496
rect 22277 3438 24000 3440
rect 22277 3435 22343 3438
rect 23200 3408 24000 3438
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 23200 2864 24000 2984
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 0 2320 800 2440
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
rect 0 1730 800 1760
rect 1577 1730 1643 1733
rect 0 1728 1643 1730
rect 0 1672 1582 1728
rect 1638 1672 1643 1728
rect 0 1670 1643 1672
rect 0 1640 800 1670
rect 1577 1667 1643 1670
rect 0 1050 800 1080
rect 1393 1050 1459 1053
rect 0 1048 1459 1050
rect 0 992 1398 1048
rect 1454 992 1459 1048
rect 0 990 1459 992
rect 0 960 800 990
rect 1393 987 1459 990
<< via3 >>
rect 3666 27772 3730 27776
rect 3666 27716 3670 27772
rect 3670 27716 3726 27772
rect 3726 27716 3730 27772
rect 3666 27712 3730 27716
rect 3746 27772 3810 27776
rect 3746 27716 3750 27772
rect 3750 27716 3806 27772
rect 3806 27716 3810 27772
rect 3746 27712 3810 27716
rect 3826 27772 3890 27776
rect 3826 27716 3830 27772
rect 3830 27716 3886 27772
rect 3886 27716 3890 27772
rect 3826 27712 3890 27716
rect 3906 27772 3970 27776
rect 3906 27716 3910 27772
rect 3910 27716 3966 27772
rect 3966 27716 3970 27772
rect 3906 27712 3970 27716
rect 9094 27772 9158 27776
rect 9094 27716 9098 27772
rect 9098 27716 9154 27772
rect 9154 27716 9158 27772
rect 9094 27712 9158 27716
rect 9174 27772 9238 27776
rect 9174 27716 9178 27772
rect 9178 27716 9234 27772
rect 9234 27716 9238 27772
rect 9174 27712 9238 27716
rect 9254 27772 9318 27776
rect 9254 27716 9258 27772
rect 9258 27716 9314 27772
rect 9314 27716 9318 27772
rect 9254 27712 9318 27716
rect 9334 27772 9398 27776
rect 9334 27716 9338 27772
rect 9338 27716 9394 27772
rect 9394 27716 9398 27772
rect 9334 27712 9398 27716
rect 14522 27772 14586 27776
rect 14522 27716 14526 27772
rect 14526 27716 14582 27772
rect 14582 27716 14586 27772
rect 14522 27712 14586 27716
rect 14602 27772 14666 27776
rect 14602 27716 14606 27772
rect 14606 27716 14662 27772
rect 14662 27716 14666 27772
rect 14602 27712 14666 27716
rect 14682 27772 14746 27776
rect 14682 27716 14686 27772
rect 14686 27716 14742 27772
rect 14742 27716 14746 27772
rect 14682 27712 14746 27716
rect 14762 27772 14826 27776
rect 14762 27716 14766 27772
rect 14766 27716 14822 27772
rect 14822 27716 14826 27772
rect 14762 27712 14826 27716
rect 19950 27772 20014 27776
rect 19950 27716 19954 27772
rect 19954 27716 20010 27772
rect 20010 27716 20014 27772
rect 19950 27712 20014 27716
rect 20030 27772 20094 27776
rect 20030 27716 20034 27772
rect 20034 27716 20090 27772
rect 20090 27716 20094 27772
rect 20030 27712 20094 27716
rect 20110 27772 20174 27776
rect 20110 27716 20114 27772
rect 20114 27716 20170 27772
rect 20170 27716 20174 27772
rect 20110 27712 20174 27716
rect 20190 27772 20254 27776
rect 20190 27716 20194 27772
rect 20194 27716 20250 27772
rect 20250 27716 20254 27772
rect 20190 27712 20254 27716
rect 6380 27228 6444 27232
rect 6380 27172 6384 27228
rect 6384 27172 6440 27228
rect 6440 27172 6444 27228
rect 6380 27168 6444 27172
rect 6460 27228 6524 27232
rect 6460 27172 6464 27228
rect 6464 27172 6520 27228
rect 6520 27172 6524 27228
rect 6460 27168 6524 27172
rect 6540 27228 6604 27232
rect 6540 27172 6544 27228
rect 6544 27172 6600 27228
rect 6600 27172 6604 27228
rect 6540 27168 6604 27172
rect 6620 27228 6684 27232
rect 6620 27172 6624 27228
rect 6624 27172 6680 27228
rect 6680 27172 6684 27228
rect 6620 27168 6684 27172
rect 11808 27228 11872 27232
rect 11808 27172 11812 27228
rect 11812 27172 11868 27228
rect 11868 27172 11872 27228
rect 11808 27168 11872 27172
rect 11888 27228 11952 27232
rect 11888 27172 11892 27228
rect 11892 27172 11948 27228
rect 11948 27172 11952 27228
rect 11888 27168 11952 27172
rect 11968 27228 12032 27232
rect 11968 27172 11972 27228
rect 11972 27172 12028 27228
rect 12028 27172 12032 27228
rect 11968 27168 12032 27172
rect 12048 27228 12112 27232
rect 12048 27172 12052 27228
rect 12052 27172 12108 27228
rect 12108 27172 12112 27228
rect 12048 27168 12112 27172
rect 17236 27228 17300 27232
rect 17236 27172 17240 27228
rect 17240 27172 17296 27228
rect 17296 27172 17300 27228
rect 17236 27168 17300 27172
rect 17316 27228 17380 27232
rect 17316 27172 17320 27228
rect 17320 27172 17376 27228
rect 17376 27172 17380 27228
rect 17316 27168 17380 27172
rect 17396 27228 17460 27232
rect 17396 27172 17400 27228
rect 17400 27172 17456 27228
rect 17456 27172 17460 27228
rect 17396 27168 17460 27172
rect 17476 27228 17540 27232
rect 17476 27172 17480 27228
rect 17480 27172 17536 27228
rect 17536 27172 17540 27228
rect 17476 27168 17540 27172
rect 22664 27228 22728 27232
rect 22664 27172 22668 27228
rect 22668 27172 22724 27228
rect 22724 27172 22728 27228
rect 22664 27168 22728 27172
rect 22744 27228 22808 27232
rect 22744 27172 22748 27228
rect 22748 27172 22804 27228
rect 22804 27172 22808 27228
rect 22744 27168 22808 27172
rect 22824 27228 22888 27232
rect 22824 27172 22828 27228
rect 22828 27172 22884 27228
rect 22884 27172 22888 27228
rect 22824 27168 22888 27172
rect 22904 27228 22968 27232
rect 22904 27172 22908 27228
rect 22908 27172 22964 27228
rect 22964 27172 22968 27228
rect 22904 27168 22968 27172
rect 3666 26684 3730 26688
rect 3666 26628 3670 26684
rect 3670 26628 3726 26684
rect 3726 26628 3730 26684
rect 3666 26624 3730 26628
rect 3746 26684 3810 26688
rect 3746 26628 3750 26684
rect 3750 26628 3806 26684
rect 3806 26628 3810 26684
rect 3746 26624 3810 26628
rect 3826 26684 3890 26688
rect 3826 26628 3830 26684
rect 3830 26628 3886 26684
rect 3886 26628 3890 26684
rect 3826 26624 3890 26628
rect 3906 26684 3970 26688
rect 3906 26628 3910 26684
rect 3910 26628 3966 26684
rect 3966 26628 3970 26684
rect 3906 26624 3970 26628
rect 9094 26684 9158 26688
rect 9094 26628 9098 26684
rect 9098 26628 9154 26684
rect 9154 26628 9158 26684
rect 9094 26624 9158 26628
rect 9174 26684 9238 26688
rect 9174 26628 9178 26684
rect 9178 26628 9234 26684
rect 9234 26628 9238 26684
rect 9174 26624 9238 26628
rect 9254 26684 9318 26688
rect 9254 26628 9258 26684
rect 9258 26628 9314 26684
rect 9314 26628 9318 26684
rect 9254 26624 9318 26628
rect 9334 26684 9398 26688
rect 9334 26628 9338 26684
rect 9338 26628 9394 26684
rect 9394 26628 9398 26684
rect 9334 26624 9398 26628
rect 14522 26684 14586 26688
rect 14522 26628 14526 26684
rect 14526 26628 14582 26684
rect 14582 26628 14586 26684
rect 14522 26624 14586 26628
rect 14602 26684 14666 26688
rect 14602 26628 14606 26684
rect 14606 26628 14662 26684
rect 14662 26628 14666 26684
rect 14602 26624 14666 26628
rect 14682 26684 14746 26688
rect 14682 26628 14686 26684
rect 14686 26628 14742 26684
rect 14742 26628 14746 26684
rect 14682 26624 14746 26628
rect 14762 26684 14826 26688
rect 14762 26628 14766 26684
rect 14766 26628 14822 26684
rect 14822 26628 14826 26684
rect 14762 26624 14826 26628
rect 19950 26684 20014 26688
rect 19950 26628 19954 26684
rect 19954 26628 20010 26684
rect 20010 26628 20014 26684
rect 19950 26624 20014 26628
rect 20030 26684 20094 26688
rect 20030 26628 20034 26684
rect 20034 26628 20090 26684
rect 20090 26628 20094 26684
rect 20030 26624 20094 26628
rect 20110 26684 20174 26688
rect 20110 26628 20114 26684
rect 20114 26628 20170 26684
rect 20170 26628 20174 26684
rect 20110 26624 20174 26628
rect 20190 26684 20254 26688
rect 20190 26628 20194 26684
rect 20194 26628 20250 26684
rect 20250 26628 20254 26684
rect 20190 26624 20254 26628
rect 21404 26420 21468 26484
rect 4108 26284 4172 26348
rect 6380 26140 6444 26144
rect 6380 26084 6384 26140
rect 6384 26084 6440 26140
rect 6440 26084 6444 26140
rect 6380 26080 6444 26084
rect 6460 26140 6524 26144
rect 6460 26084 6464 26140
rect 6464 26084 6520 26140
rect 6520 26084 6524 26140
rect 6460 26080 6524 26084
rect 6540 26140 6604 26144
rect 6540 26084 6544 26140
rect 6544 26084 6600 26140
rect 6600 26084 6604 26140
rect 6540 26080 6604 26084
rect 6620 26140 6684 26144
rect 6620 26084 6624 26140
rect 6624 26084 6680 26140
rect 6680 26084 6684 26140
rect 6620 26080 6684 26084
rect 11808 26140 11872 26144
rect 11808 26084 11812 26140
rect 11812 26084 11868 26140
rect 11868 26084 11872 26140
rect 11808 26080 11872 26084
rect 11888 26140 11952 26144
rect 11888 26084 11892 26140
rect 11892 26084 11948 26140
rect 11948 26084 11952 26140
rect 11888 26080 11952 26084
rect 11968 26140 12032 26144
rect 11968 26084 11972 26140
rect 11972 26084 12028 26140
rect 12028 26084 12032 26140
rect 11968 26080 12032 26084
rect 12048 26140 12112 26144
rect 12048 26084 12052 26140
rect 12052 26084 12108 26140
rect 12108 26084 12112 26140
rect 12048 26080 12112 26084
rect 17236 26140 17300 26144
rect 17236 26084 17240 26140
rect 17240 26084 17296 26140
rect 17296 26084 17300 26140
rect 17236 26080 17300 26084
rect 17316 26140 17380 26144
rect 17316 26084 17320 26140
rect 17320 26084 17376 26140
rect 17376 26084 17380 26140
rect 17316 26080 17380 26084
rect 17396 26140 17460 26144
rect 17396 26084 17400 26140
rect 17400 26084 17456 26140
rect 17456 26084 17460 26140
rect 17396 26080 17460 26084
rect 17476 26140 17540 26144
rect 17476 26084 17480 26140
rect 17480 26084 17536 26140
rect 17536 26084 17540 26140
rect 17476 26080 17540 26084
rect 22664 26140 22728 26144
rect 22664 26084 22668 26140
rect 22668 26084 22724 26140
rect 22724 26084 22728 26140
rect 22664 26080 22728 26084
rect 22744 26140 22808 26144
rect 22744 26084 22748 26140
rect 22748 26084 22804 26140
rect 22804 26084 22808 26140
rect 22744 26080 22808 26084
rect 22824 26140 22888 26144
rect 22824 26084 22828 26140
rect 22828 26084 22884 26140
rect 22884 26084 22888 26140
rect 22824 26080 22888 26084
rect 22904 26140 22968 26144
rect 22904 26084 22908 26140
rect 22908 26084 22964 26140
rect 22964 26084 22968 26140
rect 22904 26080 22968 26084
rect 3666 25596 3730 25600
rect 3666 25540 3670 25596
rect 3670 25540 3726 25596
rect 3726 25540 3730 25596
rect 3666 25536 3730 25540
rect 3746 25596 3810 25600
rect 3746 25540 3750 25596
rect 3750 25540 3806 25596
rect 3806 25540 3810 25596
rect 3746 25536 3810 25540
rect 3826 25596 3890 25600
rect 3826 25540 3830 25596
rect 3830 25540 3886 25596
rect 3886 25540 3890 25596
rect 3826 25536 3890 25540
rect 3906 25596 3970 25600
rect 3906 25540 3910 25596
rect 3910 25540 3966 25596
rect 3966 25540 3970 25596
rect 3906 25536 3970 25540
rect 9094 25596 9158 25600
rect 9094 25540 9098 25596
rect 9098 25540 9154 25596
rect 9154 25540 9158 25596
rect 9094 25536 9158 25540
rect 9174 25596 9238 25600
rect 9174 25540 9178 25596
rect 9178 25540 9234 25596
rect 9234 25540 9238 25596
rect 9174 25536 9238 25540
rect 9254 25596 9318 25600
rect 9254 25540 9258 25596
rect 9258 25540 9314 25596
rect 9314 25540 9318 25596
rect 9254 25536 9318 25540
rect 9334 25596 9398 25600
rect 9334 25540 9338 25596
rect 9338 25540 9394 25596
rect 9394 25540 9398 25596
rect 9334 25536 9398 25540
rect 14522 25596 14586 25600
rect 14522 25540 14526 25596
rect 14526 25540 14582 25596
rect 14582 25540 14586 25596
rect 14522 25536 14586 25540
rect 14602 25596 14666 25600
rect 14602 25540 14606 25596
rect 14606 25540 14662 25596
rect 14662 25540 14666 25596
rect 14602 25536 14666 25540
rect 14682 25596 14746 25600
rect 14682 25540 14686 25596
rect 14686 25540 14742 25596
rect 14742 25540 14746 25596
rect 14682 25536 14746 25540
rect 14762 25596 14826 25600
rect 14762 25540 14766 25596
rect 14766 25540 14822 25596
rect 14822 25540 14826 25596
rect 14762 25536 14826 25540
rect 19950 25596 20014 25600
rect 19950 25540 19954 25596
rect 19954 25540 20010 25596
rect 20010 25540 20014 25596
rect 19950 25536 20014 25540
rect 20030 25596 20094 25600
rect 20030 25540 20034 25596
rect 20034 25540 20090 25596
rect 20090 25540 20094 25596
rect 20030 25536 20094 25540
rect 20110 25596 20174 25600
rect 20110 25540 20114 25596
rect 20114 25540 20170 25596
rect 20170 25540 20174 25596
rect 20110 25536 20174 25540
rect 20190 25596 20254 25600
rect 20190 25540 20194 25596
rect 20194 25540 20250 25596
rect 20250 25540 20254 25596
rect 20190 25536 20254 25540
rect 6380 25052 6444 25056
rect 6380 24996 6384 25052
rect 6384 24996 6440 25052
rect 6440 24996 6444 25052
rect 6380 24992 6444 24996
rect 6460 25052 6524 25056
rect 6460 24996 6464 25052
rect 6464 24996 6520 25052
rect 6520 24996 6524 25052
rect 6460 24992 6524 24996
rect 6540 25052 6604 25056
rect 6540 24996 6544 25052
rect 6544 24996 6600 25052
rect 6600 24996 6604 25052
rect 6540 24992 6604 24996
rect 6620 25052 6684 25056
rect 6620 24996 6624 25052
rect 6624 24996 6680 25052
rect 6680 24996 6684 25052
rect 6620 24992 6684 24996
rect 11808 25052 11872 25056
rect 11808 24996 11812 25052
rect 11812 24996 11868 25052
rect 11868 24996 11872 25052
rect 11808 24992 11872 24996
rect 11888 25052 11952 25056
rect 11888 24996 11892 25052
rect 11892 24996 11948 25052
rect 11948 24996 11952 25052
rect 11888 24992 11952 24996
rect 11968 25052 12032 25056
rect 11968 24996 11972 25052
rect 11972 24996 12028 25052
rect 12028 24996 12032 25052
rect 11968 24992 12032 24996
rect 12048 25052 12112 25056
rect 12048 24996 12052 25052
rect 12052 24996 12108 25052
rect 12108 24996 12112 25052
rect 12048 24992 12112 24996
rect 17236 25052 17300 25056
rect 17236 24996 17240 25052
rect 17240 24996 17296 25052
rect 17296 24996 17300 25052
rect 17236 24992 17300 24996
rect 17316 25052 17380 25056
rect 17316 24996 17320 25052
rect 17320 24996 17376 25052
rect 17376 24996 17380 25052
rect 17316 24992 17380 24996
rect 17396 25052 17460 25056
rect 17396 24996 17400 25052
rect 17400 24996 17456 25052
rect 17456 24996 17460 25052
rect 17396 24992 17460 24996
rect 17476 25052 17540 25056
rect 17476 24996 17480 25052
rect 17480 24996 17536 25052
rect 17536 24996 17540 25052
rect 17476 24992 17540 24996
rect 22664 25052 22728 25056
rect 22664 24996 22668 25052
rect 22668 24996 22724 25052
rect 22724 24996 22728 25052
rect 22664 24992 22728 24996
rect 22744 25052 22808 25056
rect 22744 24996 22748 25052
rect 22748 24996 22804 25052
rect 22804 24996 22808 25052
rect 22744 24992 22808 24996
rect 22824 25052 22888 25056
rect 22824 24996 22828 25052
rect 22828 24996 22884 25052
rect 22884 24996 22888 25052
rect 22824 24992 22888 24996
rect 22904 25052 22968 25056
rect 22904 24996 22908 25052
rect 22908 24996 22964 25052
rect 22964 24996 22968 25052
rect 22904 24992 22968 24996
rect 4292 24924 4356 24988
rect 3666 24508 3730 24512
rect 3666 24452 3670 24508
rect 3670 24452 3726 24508
rect 3726 24452 3730 24508
rect 3666 24448 3730 24452
rect 3746 24508 3810 24512
rect 3746 24452 3750 24508
rect 3750 24452 3806 24508
rect 3806 24452 3810 24508
rect 3746 24448 3810 24452
rect 3826 24508 3890 24512
rect 3826 24452 3830 24508
rect 3830 24452 3886 24508
rect 3886 24452 3890 24508
rect 3826 24448 3890 24452
rect 3906 24508 3970 24512
rect 3906 24452 3910 24508
rect 3910 24452 3966 24508
rect 3966 24452 3970 24508
rect 3906 24448 3970 24452
rect 9094 24508 9158 24512
rect 9094 24452 9098 24508
rect 9098 24452 9154 24508
rect 9154 24452 9158 24508
rect 9094 24448 9158 24452
rect 9174 24508 9238 24512
rect 9174 24452 9178 24508
rect 9178 24452 9234 24508
rect 9234 24452 9238 24508
rect 9174 24448 9238 24452
rect 9254 24508 9318 24512
rect 9254 24452 9258 24508
rect 9258 24452 9314 24508
rect 9314 24452 9318 24508
rect 9254 24448 9318 24452
rect 9334 24508 9398 24512
rect 9334 24452 9338 24508
rect 9338 24452 9394 24508
rect 9394 24452 9398 24508
rect 9334 24448 9398 24452
rect 14522 24508 14586 24512
rect 14522 24452 14526 24508
rect 14526 24452 14582 24508
rect 14582 24452 14586 24508
rect 14522 24448 14586 24452
rect 14602 24508 14666 24512
rect 14602 24452 14606 24508
rect 14606 24452 14662 24508
rect 14662 24452 14666 24508
rect 14602 24448 14666 24452
rect 14682 24508 14746 24512
rect 14682 24452 14686 24508
rect 14686 24452 14742 24508
rect 14742 24452 14746 24508
rect 14682 24448 14746 24452
rect 14762 24508 14826 24512
rect 14762 24452 14766 24508
rect 14766 24452 14822 24508
rect 14822 24452 14826 24508
rect 14762 24448 14826 24452
rect 19950 24508 20014 24512
rect 19950 24452 19954 24508
rect 19954 24452 20010 24508
rect 20010 24452 20014 24508
rect 19950 24448 20014 24452
rect 20030 24508 20094 24512
rect 20030 24452 20034 24508
rect 20034 24452 20090 24508
rect 20090 24452 20094 24508
rect 20030 24448 20094 24452
rect 20110 24508 20174 24512
rect 20110 24452 20114 24508
rect 20114 24452 20170 24508
rect 20170 24452 20174 24508
rect 20110 24448 20174 24452
rect 20190 24508 20254 24512
rect 20190 24452 20194 24508
rect 20194 24452 20250 24508
rect 20250 24452 20254 24508
rect 20190 24448 20254 24452
rect 6380 23964 6444 23968
rect 6380 23908 6384 23964
rect 6384 23908 6440 23964
rect 6440 23908 6444 23964
rect 6380 23904 6444 23908
rect 6460 23964 6524 23968
rect 6460 23908 6464 23964
rect 6464 23908 6520 23964
rect 6520 23908 6524 23964
rect 6460 23904 6524 23908
rect 6540 23964 6604 23968
rect 6540 23908 6544 23964
rect 6544 23908 6600 23964
rect 6600 23908 6604 23964
rect 6540 23904 6604 23908
rect 6620 23964 6684 23968
rect 6620 23908 6624 23964
rect 6624 23908 6680 23964
rect 6680 23908 6684 23964
rect 6620 23904 6684 23908
rect 11808 23964 11872 23968
rect 11808 23908 11812 23964
rect 11812 23908 11868 23964
rect 11868 23908 11872 23964
rect 11808 23904 11872 23908
rect 11888 23964 11952 23968
rect 11888 23908 11892 23964
rect 11892 23908 11948 23964
rect 11948 23908 11952 23964
rect 11888 23904 11952 23908
rect 11968 23964 12032 23968
rect 11968 23908 11972 23964
rect 11972 23908 12028 23964
rect 12028 23908 12032 23964
rect 11968 23904 12032 23908
rect 12048 23964 12112 23968
rect 12048 23908 12052 23964
rect 12052 23908 12108 23964
rect 12108 23908 12112 23964
rect 12048 23904 12112 23908
rect 17236 23964 17300 23968
rect 17236 23908 17240 23964
rect 17240 23908 17296 23964
rect 17296 23908 17300 23964
rect 17236 23904 17300 23908
rect 17316 23964 17380 23968
rect 17316 23908 17320 23964
rect 17320 23908 17376 23964
rect 17376 23908 17380 23964
rect 17316 23904 17380 23908
rect 17396 23964 17460 23968
rect 17396 23908 17400 23964
rect 17400 23908 17456 23964
rect 17456 23908 17460 23964
rect 17396 23904 17460 23908
rect 17476 23964 17540 23968
rect 17476 23908 17480 23964
rect 17480 23908 17536 23964
rect 17536 23908 17540 23964
rect 17476 23904 17540 23908
rect 22664 23964 22728 23968
rect 22664 23908 22668 23964
rect 22668 23908 22724 23964
rect 22724 23908 22728 23964
rect 22664 23904 22728 23908
rect 22744 23964 22808 23968
rect 22744 23908 22748 23964
rect 22748 23908 22804 23964
rect 22804 23908 22808 23964
rect 22744 23904 22808 23908
rect 22824 23964 22888 23968
rect 22824 23908 22828 23964
rect 22828 23908 22884 23964
rect 22884 23908 22888 23964
rect 22824 23904 22888 23908
rect 22904 23964 22968 23968
rect 22904 23908 22908 23964
rect 22908 23908 22964 23964
rect 22964 23908 22968 23964
rect 22904 23904 22968 23908
rect 3666 23420 3730 23424
rect 3666 23364 3670 23420
rect 3670 23364 3726 23420
rect 3726 23364 3730 23420
rect 3666 23360 3730 23364
rect 3746 23420 3810 23424
rect 3746 23364 3750 23420
rect 3750 23364 3806 23420
rect 3806 23364 3810 23420
rect 3746 23360 3810 23364
rect 3826 23420 3890 23424
rect 3826 23364 3830 23420
rect 3830 23364 3886 23420
rect 3886 23364 3890 23420
rect 3826 23360 3890 23364
rect 3906 23420 3970 23424
rect 3906 23364 3910 23420
rect 3910 23364 3966 23420
rect 3966 23364 3970 23420
rect 3906 23360 3970 23364
rect 9094 23420 9158 23424
rect 9094 23364 9098 23420
rect 9098 23364 9154 23420
rect 9154 23364 9158 23420
rect 9094 23360 9158 23364
rect 9174 23420 9238 23424
rect 9174 23364 9178 23420
rect 9178 23364 9234 23420
rect 9234 23364 9238 23420
rect 9174 23360 9238 23364
rect 9254 23420 9318 23424
rect 9254 23364 9258 23420
rect 9258 23364 9314 23420
rect 9314 23364 9318 23420
rect 9254 23360 9318 23364
rect 9334 23420 9398 23424
rect 9334 23364 9338 23420
rect 9338 23364 9394 23420
rect 9394 23364 9398 23420
rect 9334 23360 9398 23364
rect 14522 23420 14586 23424
rect 14522 23364 14526 23420
rect 14526 23364 14582 23420
rect 14582 23364 14586 23420
rect 14522 23360 14586 23364
rect 14602 23420 14666 23424
rect 14602 23364 14606 23420
rect 14606 23364 14662 23420
rect 14662 23364 14666 23420
rect 14602 23360 14666 23364
rect 14682 23420 14746 23424
rect 14682 23364 14686 23420
rect 14686 23364 14742 23420
rect 14742 23364 14746 23420
rect 14682 23360 14746 23364
rect 14762 23420 14826 23424
rect 14762 23364 14766 23420
rect 14766 23364 14822 23420
rect 14822 23364 14826 23420
rect 14762 23360 14826 23364
rect 19950 23420 20014 23424
rect 19950 23364 19954 23420
rect 19954 23364 20010 23420
rect 20010 23364 20014 23420
rect 19950 23360 20014 23364
rect 20030 23420 20094 23424
rect 20030 23364 20034 23420
rect 20034 23364 20090 23420
rect 20090 23364 20094 23420
rect 20030 23360 20094 23364
rect 20110 23420 20174 23424
rect 20110 23364 20114 23420
rect 20114 23364 20170 23420
rect 20170 23364 20174 23420
rect 20110 23360 20174 23364
rect 20190 23420 20254 23424
rect 20190 23364 20194 23420
rect 20194 23364 20250 23420
rect 20250 23364 20254 23420
rect 20190 23360 20254 23364
rect 4108 23216 4172 23220
rect 4108 23160 4158 23216
rect 4158 23160 4172 23216
rect 4108 23156 4172 23160
rect 6380 22876 6444 22880
rect 6380 22820 6384 22876
rect 6384 22820 6440 22876
rect 6440 22820 6444 22876
rect 6380 22816 6444 22820
rect 6460 22876 6524 22880
rect 6460 22820 6464 22876
rect 6464 22820 6520 22876
rect 6520 22820 6524 22876
rect 6460 22816 6524 22820
rect 6540 22876 6604 22880
rect 6540 22820 6544 22876
rect 6544 22820 6600 22876
rect 6600 22820 6604 22876
rect 6540 22816 6604 22820
rect 6620 22876 6684 22880
rect 6620 22820 6624 22876
rect 6624 22820 6680 22876
rect 6680 22820 6684 22876
rect 6620 22816 6684 22820
rect 11808 22876 11872 22880
rect 11808 22820 11812 22876
rect 11812 22820 11868 22876
rect 11868 22820 11872 22876
rect 11808 22816 11872 22820
rect 11888 22876 11952 22880
rect 11888 22820 11892 22876
rect 11892 22820 11948 22876
rect 11948 22820 11952 22876
rect 11888 22816 11952 22820
rect 11968 22876 12032 22880
rect 11968 22820 11972 22876
rect 11972 22820 12028 22876
rect 12028 22820 12032 22876
rect 11968 22816 12032 22820
rect 12048 22876 12112 22880
rect 12048 22820 12052 22876
rect 12052 22820 12108 22876
rect 12108 22820 12112 22876
rect 12048 22816 12112 22820
rect 17236 22876 17300 22880
rect 17236 22820 17240 22876
rect 17240 22820 17296 22876
rect 17296 22820 17300 22876
rect 17236 22816 17300 22820
rect 17316 22876 17380 22880
rect 17316 22820 17320 22876
rect 17320 22820 17376 22876
rect 17376 22820 17380 22876
rect 17316 22816 17380 22820
rect 17396 22876 17460 22880
rect 17396 22820 17400 22876
rect 17400 22820 17456 22876
rect 17456 22820 17460 22876
rect 17396 22816 17460 22820
rect 17476 22876 17540 22880
rect 17476 22820 17480 22876
rect 17480 22820 17536 22876
rect 17536 22820 17540 22876
rect 17476 22816 17540 22820
rect 22664 22876 22728 22880
rect 22664 22820 22668 22876
rect 22668 22820 22724 22876
rect 22724 22820 22728 22876
rect 22664 22816 22728 22820
rect 22744 22876 22808 22880
rect 22744 22820 22748 22876
rect 22748 22820 22804 22876
rect 22804 22820 22808 22876
rect 22744 22816 22808 22820
rect 22824 22876 22888 22880
rect 22824 22820 22828 22876
rect 22828 22820 22884 22876
rect 22884 22820 22888 22876
rect 22824 22816 22888 22820
rect 22904 22876 22968 22880
rect 22904 22820 22908 22876
rect 22908 22820 22964 22876
rect 22964 22820 22968 22876
rect 22904 22816 22968 22820
rect 3666 22332 3730 22336
rect 3666 22276 3670 22332
rect 3670 22276 3726 22332
rect 3726 22276 3730 22332
rect 3666 22272 3730 22276
rect 3746 22332 3810 22336
rect 3746 22276 3750 22332
rect 3750 22276 3806 22332
rect 3806 22276 3810 22332
rect 3746 22272 3810 22276
rect 3826 22332 3890 22336
rect 3826 22276 3830 22332
rect 3830 22276 3886 22332
rect 3886 22276 3890 22332
rect 3826 22272 3890 22276
rect 3906 22332 3970 22336
rect 3906 22276 3910 22332
rect 3910 22276 3966 22332
rect 3966 22276 3970 22332
rect 3906 22272 3970 22276
rect 9094 22332 9158 22336
rect 9094 22276 9098 22332
rect 9098 22276 9154 22332
rect 9154 22276 9158 22332
rect 9094 22272 9158 22276
rect 9174 22332 9238 22336
rect 9174 22276 9178 22332
rect 9178 22276 9234 22332
rect 9234 22276 9238 22332
rect 9174 22272 9238 22276
rect 9254 22332 9318 22336
rect 9254 22276 9258 22332
rect 9258 22276 9314 22332
rect 9314 22276 9318 22332
rect 9254 22272 9318 22276
rect 9334 22332 9398 22336
rect 9334 22276 9338 22332
rect 9338 22276 9394 22332
rect 9394 22276 9398 22332
rect 9334 22272 9398 22276
rect 14522 22332 14586 22336
rect 14522 22276 14526 22332
rect 14526 22276 14582 22332
rect 14582 22276 14586 22332
rect 14522 22272 14586 22276
rect 14602 22332 14666 22336
rect 14602 22276 14606 22332
rect 14606 22276 14662 22332
rect 14662 22276 14666 22332
rect 14602 22272 14666 22276
rect 14682 22332 14746 22336
rect 14682 22276 14686 22332
rect 14686 22276 14742 22332
rect 14742 22276 14746 22332
rect 14682 22272 14746 22276
rect 14762 22332 14826 22336
rect 14762 22276 14766 22332
rect 14766 22276 14822 22332
rect 14822 22276 14826 22332
rect 14762 22272 14826 22276
rect 19950 22332 20014 22336
rect 19950 22276 19954 22332
rect 19954 22276 20010 22332
rect 20010 22276 20014 22332
rect 19950 22272 20014 22276
rect 20030 22332 20094 22336
rect 20030 22276 20034 22332
rect 20034 22276 20090 22332
rect 20090 22276 20094 22332
rect 20030 22272 20094 22276
rect 20110 22332 20174 22336
rect 20110 22276 20114 22332
rect 20114 22276 20170 22332
rect 20170 22276 20174 22332
rect 20110 22272 20174 22276
rect 20190 22332 20254 22336
rect 20190 22276 20194 22332
rect 20194 22276 20250 22332
rect 20250 22276 20254 22332
rect 20190 22272 20254 22276
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 4292 21660 4356 21724
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 21404 20572 21468 20636
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 5028 19348 5092 19412
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 4292 18124 4356 18188
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 5028 15736 5092 15740
rect 5028 15680 5078 15736
rect 5078 15680 5092 15736
rect 5028 15676 5092 15680
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 4292 14512 4356 14516
rect 4292 14456 4342 14512
rect 4342 14456 4356 14512
rect 4292 14452 4356 14456
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 27776 3978 27792
rect 3658 27712 3666 27776
rect 3730 27712 3746 27776
rect 3810 27712 3826 27776
rect 3890 27712 3906 27776
rect 3970 27712 3978 27776
rect 3658 26688 3978 27712
rect 3658 26624 3666 26688
rect 3730 26624 3746 26688
rect 3810 26624 3826 26688
rect 3890 26624 3906 26688
rect 3970 26624 3978 26688
rect 3658 25600 3978 26624
rect 6372 27232 6692 27792
rect 6372 27168 6380 27232
rect 6444 27168 6460 27232
rect 6524 27168 6540 27232
rect 6604 27168 6620 27232
rect 6684 27168 6692 27232
rect 4107 26348 4173 26349
rect 4107 26284 4108 26348
rect 4172 26284 4173 26348
rect 4107 26283 4173 26284
rect 3658 25536 3666 25600
rect 3730 25536 3746 25600
rect 3810 25536 3826 25600
rect 3890 25536 3906 25600
rect 3970 25536 3978 25600
rect 3658 24512 3978 25536
rect 3658 24448 3666 24512
rect 3730 24448 3746 24512
rect 3810 24448 3826 24512
rect 3890 24448 3906 24512
rect 3970 24448 3978 24512
rect 3658 23424 3978 24448
rect 3658 23360 3666 23424
rect 3730 23360 3746 23424
rect 3810 23360 3826 23424
rect 3890 23360 3906 23424
rect 3970 23360 3978 23424
rect 3658 22336 3978 23360
rect 4110 23221 4170 26283
rect 6372 26144 6692 27168
rect 6372 26080 6380 26144
rect 6444 26080 6460 26144
rect 6524 26080 6540 26144
rect 6604 26080 6620 26144
rect 6684 26080 6692 26144
rect 6372 25056 6692 26080
rect 6372 24992 6380 25056
rect 6444 24992 6460 25056
rect 6524 24992 6540 25056
rect 6604 24992 6620 25056
rect 6684 24992 6692 25056
rect 4291 24988 4357 24989
rect 4291 24924 4292 24988
rect 4356 24924 4357 24988
rect 4291 24923 4357 24924
rect 4107 23220 4173 23221
rect 4107 23156 4108 23220
rect 4172 23156 4173 23220
rect 4107 23155 4173 23156
rect 3658 22272 3666 22336
rect 3730 22272 3746 22336
rect 3810 22272 3826 22336
rect 3890 22272 3906 22336
rect 3970 22272 3978 22336
rect 3658 21248 3978 22272
rect 4294 21725 4354 24923
rect 6372 23968 6692 24992
rect 6372 23904 6380 23968
rect 6444 23904 6460 23968
rect 6524 23904 6540 23968
rect 6604 23904 6620 23968
rect 6684 23904 6692 23968
rect 6372 22880 6692 23904
rect 6372 22816 6380 22880
rect 6444 22816 6460 22880
rect 6524 22816 6540 22880
rect 6604 22816 6620 22880
rect 6684 22816 6692 22880
rect 6372 21792 6692 22816
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 4291 21724 4357 21725
rect 4291 21660 4292 21724
rect 4356 21660 4357 21724
rect 4291 21659 4357 21660
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 5027 19412 5093 19413
rect 5027 19348 5028 19412
rect 5092 19348 5093 19412
rect 5027 19347 5093 19348
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 4291 18188 4357 18189
rect 4291 18124 4292 18188
rect 4356 18124 4357 18188
rect 4291 18123 4357 18124
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 4294 14517 4354 18123
rect 5030 15741 5090 19347
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 5027 15740 5093 15741
rect 5027 15676 5028 15740
rect 5092 15676 5093 15740
rect 5027 15675 5093 15676
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 4291 14516 4357 14517
rect 4291 14452 4292 14516
rect 4356 14452 4357 14516
rect 4291 14451 4357 14452
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 27776 9406 27792
rect 9086 27712 9094 27776
rect 9158 27712 9174 27776
rect 9238 27712 9254 27776
rect 9318 27712 9334 27776
rect 9398 27712 9406 27776
rect 9086 26688 9406 27712
rect 9086 26624 9094 26688
rect 9158 26624 9174 26688
rect 9238 26624 9254 26688
rect 9318 26624 9334 26688
rect 9398 26624 9406 26688
rect 9086 25600 9406 26624
rect 9086 25536 9094 25600
rect 9158 25536 9174 25600
rect 9238 25536 9254 25600
rect 9318 25536 9334 25600
rect 9398 25536 9406 25600
rect 9086 24512 9406 25536
rect 9086 24448 9094 24512
rect 9158 24448 9174 24512
rect 9238 24448 9254 24512
rect 9318 24448 9334 24512
rect 9398 24448 9406 24512
rect 9086 23424 9406 24448
rect 9086 23360 9094 23424
rect 9158 23360 9174 23424
rect 9238 23360 9254 23424
rect 9318 23360 9334 23424
rect 9398 23360 9406 23424
rect 9086 22336 9406 23360
rect 9086 22272 9094 22336
rect 9158 22272 9174 22336
rect 9238 22272 9254 22336
rect 9318 22272 9334 22336
rect 9398 22272 9406 22336
rect 9086 21248 9406 22272
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 27232 12120 27792
rect 11800 27168 11808 27232
rect 11872 27168 11888 27232
rect 11952 27168 11968 27232
rect 12032 27168 12048 27232
rect 12112 27168 12120 27232
rect 11800 26144 12120 27168
rect 11800 26080 11808 26144
rect 11872 26080 11888 26144
rect 11952 26080 11968 26144
rect 12032 26080 12048 26144
rect 12112 26080 12120 26144
rect 11800 25056 12120 26080
rect 11800 24992 11808 25056
rect 11872 24992 11888 25056
rect 11952 24992 11968 25056
rect 12032 24992 12048 25056
rect 12112 24992 12120 25056
rect 11800 23968 12120 24992
rect 11800 23904 11808 23968
rect 11872 23904 11888 23968
rect 11952 23904 11968 23968
rect 12032 23904 12048 23968
rect 12112 23904 12120 23968
rect 11800 22880 12120 23904
rect 11800 22816 11808 22880
rect 11872 22816 11888 22880
rect 11952 22816 11968 22880
rect 12032 22816 12048 22880
rect 12112 22816 12120 22880
rect 11800 21792 12120 22816
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 27776 14834 27792
rect 14514 27712 14522 27776
rect 14586 27712 14602 27776
rect 14666 27712 14682 27776
rect 14746 27712 14762 27776
rect 14826 27712 14834 27776
rect 14514 26688 14834 27712
rect 14514 26624 14522 26688
rect 14586 26624 14602 26688
rect 14666 26624 14682 26688
rect 14746 26624 14762 26688
rect 14826 26624 14834 26688
rect 14514 25600 14834 26624
rect 14514 25536 14522 25600
rect 14586 25536 14602 25600
rect 14666 25536 14682 25600
rect 14746 25536 14762 25600
rect 14826 25536 14834 25600
rect 14514 24512 14834 25536
rect 14514 24448 14522 24512
rect 14586 24448 14602 24512
rect 14666 24448 14682 24512
rect 14746 24448 14762 24512
rect 14826 24448 14834 24512
rect 14514 23424 14834 24448
rect 14514 23360 14522 23424
rect 14586 23360 14602 23424
rect 14666 23360 14682 23424
rect 14746 23360 14762 23424
rect 14826 23360 14834 23424
rect 14514 22336 14834 23360
rect 14514 22272 14522 22336
rect 14586 22272 14602 22336
rect 14666 22272 14682 22336
rect 14746 22272 14762 22336
rect 14826 22272 14834 22336
rect 14514 21248 14834 22272
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 27232 17548 27792
rect 17228 27168 17236 27232
rect 17300 27168 17316 27232
rect 17380 27168 17396 27232
rect 17460 27168 17476 27232
rect 17540 27168 17548 27232
rect 17228 26144 17548 27168
rect 17228 26080 17236 26144
rect 17300 26080 17316 26144
rect 17380 26080 17396 26144
rect 17460 26080 17476 26144
rect 17540 26080 17548 26144
rect 17228 25056 17548 26080
rect 17228 24992 17236 25056
rect 17300 24992 17316 25056
rect 17380 24992 17396 25056
rect 17460 24992 17476 25056
rect 17540 24992 17548 25056
rect 17228 23968 17548 24992
rect 17228 23904 17236 23968
rect 17300 23904 17316 23968
rect 17380 23904 17396 23968
rect 17460 23904 17476 23968
rect 17540 23904 17548 23968
rect 17228 22880 17548 23904
rect 17228 22816 17236 22880
rect 17300 22816 17316 22880
rect 17380 22816 17396 22880
rect 17460 22816 17476 22880
rect 17540 22816 17548 22880
rect 17228 21792 17548 22816
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 27776 20262 27792
rect 19942 27712 19950 27776
rect 20014 27712 20030 27776
rect 20094 27712 20110 27776
rect 20174 27712 20190 27776
rect 20254 27712 20262 27776
rect 19942 26688 20262 27712
rect 19942 26624 19950 26688
rect 20014 26624 20030 26688
rect 20094 26624 20110 26688
rect 20174 26624 20190 26688
rect 20254 26624 20262 26688
rect 19942 25600 20262 26624
rect 22656 27232 22976 27792
rect 22656 27168 22664 27232
rect 22728 27168 22744 27232
rect 22808 27168 22824 27232
rect 22888 27168 22904 27232
rect 22968 27168 22976 27232
rect 21403 26484 21469 26485
rect 21403 26420 21404 26484
rect 21468 26420 21469 26484
rect 21403 26419 21469 26420
rect 19942 25536 19950 25600
rect 20014 25536 20030 25600
rect 20094 25536 20110 25600
rect 20174 25536 20190 25600
rect 20254 25536 20262 25600
rect 19942 24512 20262 25536
rect 19942 24448 19950 24512
rect 20014 24448 20030 24512
rect 20094 24448 20110 24512
rect 20174 24448 20190 24512
rect 20254 24448 20262 24512
rect 19942 23424 20262 24448
rect 19942 23360 19950 23424
rect 20014 23360 20030 23424
rect 20094 23360 20110 23424
rect 20174 23360 20190 23424
rect 20254 23360 20262 23424
rect 19942 22336 20262 23360
rect 19942 22272 19950 22336
rect 20014 22272 20030 22336
rect 20094 22272 20110 22336
rect 20174 22272 20190 22336
rect 20254 22272 20262 22336
rect 19942 21248 20262 22272
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 21406 20637 21466 26419
rect 22656 26144 22976 27168
rect 22656 26080 22664 26144
rect 22728 26080 22744 26144
rect 22808 26080 22824 26144
rect 22888 26080 22904 26144
rect 22968 26080 22976 26144
rect 22656 25056 22976 26080
rect 22656 24992 22664 25056
rect 22728 24992 22744 25056
rect 22808 24992 22824 25056
rect 22888 24992 22904 25056
rect 22968 24992 22976 25056
rect 22656 23968 22976 24992
rect 22656 23904 22664 23968
rect 22728 23904 22744 23968
rect 22808 23904 22824 23968
rect 22888 23904 22904 23968
rect 22968 23904 22976 23968
rect 22656 22880 22976 23904
rect 22656 22816 22664 22880
rect 22728 22816 22744 22880
rect 22808 22816 22824 22880
rect 22888 22816 22904 22880
rect 22968 22816 22976 22880
rect 22656 21792 22976 22816
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 21403 20636 21469 20637
rect 21403 20572 21404 20636
rect 21468 20572 21469 20636
rect 21403 20571 21469 20572
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__307__CLK pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__CLK
timestamp 1666464484
transform 1 0 5336 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__CLK
timestamp 1666464484
transform 1 0 4784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__CLK
timestamp 1666464484
transform 1 0 8004 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__CLK
timestamp 1666464484
transform -1 0 4140 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__CLK
timestamp 1666464484
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__CLK
timestamp 1666464484
transform 1 0 5428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__CLK
timestamp 1666464484
transform -1 0 4692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__CLK
timestamp 1666464484
transform -1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__CLK
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__CLK
timestamp 1666464484
transform 1 0 12328 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__CLK
timestamp 1666464484
transform 1 0 17848 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__CLK
timestamp 1666464484
transform 1 0 17388 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__CLK
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__CLK
timestamp 1666464484
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__CLK
timestamp 1666464484
transform 1 0 17664 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__CLK
timestamp 1666464484
transform -1 0 21712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__CLK
timestamp 1666464484
transform 1 0 18768 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout30_A
timestamp 1666464484
transform 1 0 9844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout31_A
timestamp 1666464484
transform 1 0 7728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 20792 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 16836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 18768 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 18216 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 20884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 16560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 15272 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 4140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 6164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 8096 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 7360 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 3864 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 3036 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1666464484
transform -1 0 4784 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1666464484
transform -1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1666464484
transform -1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1666464484
transform -1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1666464484
transform -1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1666464484
transform -1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1666464484
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1666464484
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_231
timestamp 1666464484
transform 1 0 22356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1666464484
transform 1 0 22356 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_227
timestamp 1666464484
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_231
timestamp 1666464484
transform 1 0 22356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_9
timestamp 1666464484
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_21
timestamp 1666464484
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 1666464484
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_45
timestamp 1666464484
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1666464484
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1666464484
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1666464484
transform 1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_231
timestamp 1666464484
transform 1 0 22356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 1666464484
transform 1 0 22356 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1666464484
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_14
timestamp 1666464484
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1666464484
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_231
timestamp 1666464484
transform 1 0 22356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_227
timestamp 1666464484
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1666464484
transform 1 0 22356 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1666464484
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_14
timestamp 1666464484
transform 1 0 2392 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_26
timestamp 1666464484
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_38
timestamp 1666464484
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1666464484
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 1666464484
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_8
timestamp 1666464484
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1666464484
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_22
timestamp 1666464484
transform 1 0 3128 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_34
timestamp 1666464484
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1666464484
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1666464484
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1666464484
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_227
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1666464484
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_10
timestamp 1666464484
transform 1 0 2024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1666464484
transform 1 0 2668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1666464484
transform 1 0 3312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1666464484
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1666464484
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1666464484
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1666464484
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1666464484
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1666464484
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_40
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_52
timestamp 1666464484
transform 1 0 5888 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_64
timestamp 1666464484
transform 1 0 6992 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1666464484
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1666464484
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_231
timestamp 1666464484
transform 1 0 22356 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_12
timestamp 1666464484
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1666464484
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1666464484
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_231
timestamp 1666464484
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_36
timestamp 1666464484
transform 1 0 4416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1666464484
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_52
timestamp 1666464484
transform 1 0 5888 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_64
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1666464484
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1666464484
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp 1666464484
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1666464484
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_231
timestamp 1666464484
transform 1 0 22356 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1666464484
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_39
timestamp 1666464484
transform 1 0 4692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1666464484
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1666464484
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1666464484
transform 1 0 6808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1666464484
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_72
timestamp 1666464484
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_227
timestamp 1666464484
transform 1 0 21988 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_231
timestamp 1666464484
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1666464484
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1666464484
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_64
timestamp 1666464484
transform 1 0 6992 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_76
timestamp 1666464484
transform 1 0 8096 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_88
timestamp 1666464484
transform 1 0 9200 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_100
timestamp 1666464484
transform 1 0 10304 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1666464484
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_231
timestamp 1666464484
transform 1 0 22356 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1666464484
transform 1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1666464484
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_56
timestamp 1666464484
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_63
timestamp 1666464484
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1666464484
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_227
timestamp 1666464484
transform 1 0 21988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1666464484
transform 1 0 22356 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1666464484
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_31
timestamp 1666464484
transform 1 0 3956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1666464484
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1666464484
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1666464484
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1666464484
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1666464484
transform 1 0 4416 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_43
timestamp 1666464484
transform 1 0 5060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_55
timestamp 1666464484
transform 1 0 6164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_67
timestamp 1666464484
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1666464484
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1666464484
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_231
timestamp 1666464484
transform 1 0 22356 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_12
timestamp 1666464484
transform 1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_22
timestamp 1666464484
transform 1 0 3128 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_29
timestamp 1666464484
transform 1 0 3772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_41
timestamp 1666464484
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1666464484
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_89
timestamp 1666464484
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1666464484
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1666464484
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1666464484
transform 1 0 22356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_18
timestamp 1666464484
transform 1 0 2760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1666464484
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1666464484
transform 1 0 6716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_69
timestamp 1666464484
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1666464484
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_224
timestamp 1666464484
transform 1 0 21712 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1666464484
transform 1 0 22356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_8
timestamp 1666464484
transform 1 0 1840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1666464484
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1666464484
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1666464484
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1666464484
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1666464484
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_136
timestamp 1666464484
transform 1 0 13616 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_148
timestamp 1666464484
transform 1 0 14720 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1666464484
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1666464484
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_231
timestamp 1666464484
transform 1 0 22356 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_8
timestamp 1666464484
transform 1 0 1840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1666464484
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_145
timestamp 1666464484
transform 1 0 14444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_157
timestamp 1666464484
transform 1 0 15548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_169
timestamp 1666464484
transform 1 0 16652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_181
timestamp 1666464484
transform 1 0 17756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1666464484
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1666464484
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1666464484
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_10
timestamp 1666464484
transform 1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_17
timestamp 1666464484
transform 1 0 2668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1666464484
transform 1 0 3312 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_30
timestamp 1666464484
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_42
timestamp 1666464484
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1666464484
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_84
timestamp 1666464484
transform 1 0 8832 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_96
timestamp 1666464484
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1666464484
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1666464484
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1666464484
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1666464484
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1666464484
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1666464484
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1666464484
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1666464484
transform 1 0 22356 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_12
timestamp 1666464484
transform 1 0 2208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1666464484
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 1666464484
transform 1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_39
timestamp 1666464484
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1666464484
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_66
timestamp 1666464484
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1666464484
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_116
timestamp 1666464484
transform 1 0 11776 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1666464484
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_202
timestamp 1666464484
transform 1 0 19688 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1666464484
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_231
timestamp 1666464484
transform 1 0 22356 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1666464484
transform 1 0 2208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_22
timestamp 1666464484
transform 1 0 3128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_29
timestamp 1666464484
transform 1 0 3772 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_36
timestamp 1666464484
transform 1 0 4416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_42
timestamp 1666464484
transform 1 0 4968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1666464484
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1666464484
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1666464484
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1666464484
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1666464484
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_231
timestamp 1666464484
transform 1 0 22356 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1666464484
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_36
timestamp 1666464484
transform 1 0 4416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_43
timestamp 1666464484
transform 1 0 5060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_49
timestamp 1666464484
transform 1 0 5612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_55
timestamp 1666464484
transform 1 0 6164 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1666464484
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1666464484
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1666464484
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_107
timestamp 1666464484
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_119
timestamp 1666464484
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1666464484
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_181
timestamp 1666464484
transform 1 0 17756 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_184
timestamp 1666464484
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 1666464484
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1666464484
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_231
timestamp 1666464484
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1666464484
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_41
timestamp 1666464484
transform 1 0 4876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1666464484
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1666464484
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_61
timestamp 1666464484
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_67
timestamp 1666464484
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_79
timestamp 1666464484
transform 1 0 8372 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_91
timestamp 1666464484
transform 1 0 9476 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_103
timestamp 1666464484
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1666464484
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1666464484
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1666464484
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_231
timestamp 1666464484
transform 1 0 22356 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1666464484
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_39
timestamp 1666464484
transform 1 0 4692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_48
timestamp 1666464484
transform 1 0 5520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_55
timestamp 1666464484
transform 1 0 6164 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1666464484
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1666464484
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1666464484
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1666464484
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1666464484
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1666464484
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_231
timestamp 1666464484
transform 1 0 22356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_26
timestamp 1666464484
transform 1 0 3496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_46
timestamp 1666464484
transform 1 0 5336 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1666464484
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_64
timestamp 1666464484
transform 1 0 6992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_71
timestamp 1666464484
transform 1 0 7636 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_77
timestamp 1666464484
transform 1 0 8188 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_89
timestamp 1666464484
transform 1 0 9292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_101
timestamp 1666464484
transform 1 0 10396 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1666464484
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1666464484
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1666464484
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1666464484
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1666464484
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_230
timestamp 1666464484
transform 1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1666464484
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_38
timestamp 1666464484
transform 1 0 4600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_47
timestamp 1666464484
transform 1 0 5428 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_56
timestamp 1666464484
transform 1 0 6256 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_63
timestamp 1666464484
transform 1 0 6900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1666464484
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_76
timestamp 1666464484
transform 1 0 8096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1666464484
transform 1 0 9476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_95
timestamp 1666464484
transform 1 0 9844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_102
timestamp 1666464484
transform 1 0 10488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_111
timestamp 1666464484
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1666464484
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_124
timestamp 1666464484
transform 1 0 12512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1666464484
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_171
timestamp 1666464484
transform 1 0 16836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1666464484
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1666464484
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1666464484
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_211
timestamp 1666464484
transform 1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_231
timestamp 1666464484
transform 1 0 22356 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_21
timestamp 1666464484
transform 1 0 3036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1666464484
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_42
timestamp 1666464484
transform 1 0 4968 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1666464484
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1666464484
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1666464484
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1666464484
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1666464484
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1666464484
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1666464484
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_128
timestamp 1666464484
transform 1 0 12880 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_140
timestamp 1666464484
transform 1 0 13984 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_152
timestamp 1666464484
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1666464484
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1666464484
transform 1 0 17572 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_186
timestamp 1666464484
transform 1 0 18216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1666464484
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_230
timestamp 1666464484
transform 1 0 22264 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1666464484
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_37
timestamp 1666464484
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_44
timestamp 1666464484
transform 1 0 5152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_51
timestamp 1666464484
transform 1 0 5796 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_71
timestamp 1666464484
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1666464484
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1666464484
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1666464484
transform 1 0 9476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_117
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_127
timestamp 1666464484
transform 1 0 12788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1666464484
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1666464484
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_188
timestamp 1666464484
transform 1 0 18400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1666464484
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_211
timestamp 1666464484
transform 1 0 20516 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_231
timestamp 1666464484
transform 1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_12
timestamp 1666464484
transform 1 0 2208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_22
timestamp 1666464484
transform 1 0 3128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_31
timestamp 1666464484
transform 1 0 3956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_38
timestamp 1666464484
transform 1 0 4600 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_45
timestamp 1666464484
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1666464484
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_62
timestamp 1666464484
transform 1 0 6808 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_68
timestamp 1666464484
transform 1 0 7360 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_72
timestamp 1666464484
transform 1 0 7728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_90
timestamp 1666464484
transform 1 0 9384 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1666464484
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1666464484
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1666464484
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_141
timestamp 1666464484
transform 1 0 14076 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1666464484
transform 1 0 14720 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_154
timestamp 1666464484
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_189
timestamp 1666464484
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_192
timestamp 1666464484
transform 1 0 18768 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_199
timestamp 1666464484
transform 1 0 19412 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_206
timestamp 1666464484
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1666464484
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_230
timestamp 1666464484
transform 1 0 22264 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1666464484
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_34
timestamp 1666464484
transform 1 0 4232 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_50
timestamp 1666464484
transform 1 0 5704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_57
timestamp 1666464484
transform 1 0 6348 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_64
timestamp 1666464484
transform 1 0 6992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_73
timestamp 1666464484
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1666464484
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_89
timestamp 1666464484
transform 1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1666464484
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1666464484
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1666464484
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1666464484
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1666464484
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_162
timestamp 1666464484
transform 1 0 16008 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_168
timestamp 1666464484
transform 1 0 16560 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1666464484
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_186
timestamp 1666464484
transform 1 0 18216 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_190
timestamp 1666464484
transform 1 0 18584 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1666464484
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1666464484
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1666464484
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1666464484
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_232
timestamp 1666464484
transform 1 0 22448 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_10
timestamp 1666464484
transform 1 0 2024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_17
timestamp 1666464484
transform 1 0 2668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1666464484
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_28
timestamp 1666464484
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_32
timestamp 1666464484
transform 1 0 4048 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_36
timestamp 1666464484
transform 1 0 4416 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1666464484
transform 1 0 4784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_47
timestamp 1666464484
transform 1 0 5428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1666464484
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1666464484
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1666464484
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_90
timestamp 1666464484
transform 1 0 9384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1666464484
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_142
timestamp 1666464484
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1666464484
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_160
timestamp 1666464484
transform 1 0 15824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_174
timestamp 1666464484
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_180
timestamp 1666464484
transform 1 0 17664 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1666464484
transform 1 0 18032 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1666464484
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1666464484
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_212
timestamp 1666464484
transform 1 0 20608 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_218
timestamp 1666464484
transform 1 0 21160 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_230
timestamp 1666464484
transform 1 0 22264 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_8
timestamp 1666464484
transform 1 0 1840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1666464484
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_33
timestamp 1666464484
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_40
timestamp 1666464484
transform 1 0 4784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1666464484
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_54
timestamp 1666464484
transform 1 0 6072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_57
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1666464484
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1666464484
transform 1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1666464484
transform 1 0 11224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1666464484
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1666464484
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1666464484
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_161
timestamp 1666464484
transform 1 0 15916 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 1666464484
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1666464484
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1666464484
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_181
timestamp 1666464484
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_188
timestamp 1666464484
transform 1 0 18400 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1666464484
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1666464484
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_222
timestamp 1666464484
transform 1 0 21528 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_225
timestamp 1666464484
transform 1 0 21804 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_231
timestamp 1666464484
transform 1 0 22356 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 22816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 22816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 22816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 22816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 22816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 22816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 22816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 22816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _153_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1666464484
transform 1 0 2852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _155_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1666464484
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _157_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2116 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _158_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _159_
timestamp 1666464484
transform -1 0 5796 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _160_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _162_
timestamp 1666464484
transform -1 0 3220 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _163_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _164_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4324 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _165_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _166_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _167_
timestamp 1666464484
transform 1 0 4416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _168_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _169_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _170_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6900 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _171_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5520 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1666464484
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1666464484
transform -1 0 6256 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 1666464484
transform 1 0 2576 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _175_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1666464484
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _177_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _178_
timestamp 1666464484
transform 1 0 3956 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _179_
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1666464484
transform 1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _182_
timestamp 1666464484
transform 1 0 3956 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _183_
timestamp 1666464484
transform 1 0 1564 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1666464484
transform 1 0 3128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _185_
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _186_
timestamp 1666464484
transform 1 0 2392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _187_
timestamp 1666464484
transform -1 0 5244 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _189_
timestamp 1666464484
transform -1 0 6992 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1666464484
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _191_
timestamp 1666464484
transform 1 0 1564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1666464484
transform -1 0 2668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _193_
timestamp 1666464484
transform -1 0 3956 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _194_
timestamp 1666464484
transform -1 0 4600 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _195_
timestamp 1666464484
transform -1 0 3036 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1666464484
transform -1 0 1840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 1666464484
transform 1 0 1564 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _198_
timestamp 1666464484
transform -1 0 3128 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _199_
timestamp 1666464484
transform 1 0 3404 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1666464484
transform -1 0 4416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 1666464484
transform -1 0 6992 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _202_
timestamp 1666464484
transform -1 0 2024 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _203_
timestamp 1666464484
transform 1 0 1564 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1666464484
transform 1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 1666464484
transform -1 0 5428 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 1666464484
transform -1 0 6256 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _207_
timestamp 1666464484
transform 1 0 1564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _209_
timestamp 1666464484
transform -1 0 5520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1666464484
transform -1 0 7636 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1666464484
transform 1 0 4416 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1666464484
transform 1 0 6532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _213_
timestamp 1666464484
transform 1 0 3956 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1666464484
transform 1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _215_
timestamp 1666464484
transform 1 0 11684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1666464484
transform 1 0 16836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _217_
timestamp 1666464484
transform -1 0 14076 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1666464484
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _219_
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1666464484
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _221_
timestamp 1666464484
transform -1 0 14720 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform -1 0 8372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _223_
timestamp 1666464484
transform 1 0 8740 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1666464484
transform -1 0 10488 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _225_
timestamp 1666464484
transform 1 0 8096 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 1666464484
transform -1 0 11316 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _227_
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _229_
timestamp 1666464484
transform -1 0 9384 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _230_
timestamp 1666464484
transform 1 0 9568 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _231_
timestamp 1666464484
transform -1 0 11224 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1666464484
transform -1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _233_
timestamp 1666464484
transform -1 0 7820 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _234_
timestamp 1666464484
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _235_
timestamp 1666464484
transform -1 0 7452 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1666464484
transform -1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp 1666464484
transform -1 0 10212 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1666464484
transform -1 0 6992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_
timestamp 1666464484
transform 1 0 18400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1666464484
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _241_
timestamp 1666464484
transform -1 0 22080 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1666464484
transform 1 0 17480 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _243_
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1666464484
transform -1 0 22264 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _245_
timestamp 1666464484
transform -1 0 20516 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _246_
timestamp 1666464484
transform -1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _247_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1666464484
transform -1 0 20700 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1666464484
transform 1 0 19228 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _251_
timestamp 1666464484
transform -1 0 20516 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _253_
timestamp 1666464484
transform -1 0 20516 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _254_
timestamp 1666464484
transform -1 0 21252 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _255_
timestamp 1666464484
transform 1 0 19872 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1666464484
transform -1 0 20056 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _257_
timestamp 1666464484
transform 1 0 17204 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1666464484
transform 1 0 17848 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _259_
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform -1 0 19688 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _261_
timestamp 1666464484
transform 1 0 16652 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _263_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13616 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1666464484
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1666464484
transform 1 0 21252 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1666464484
transform 1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _267_
timestamp 1666464484
transform -1 0 19688 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1666464484
transform 1 0 18584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _269_
timestamp 1666464484
transform 1 0 21804 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _270_
timestamp 1666464484
transform 1 0 19872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _271_
timestamp 1666464484
transform 1 0 17480 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1666464484
transform -1 0 21528 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1666464484
transform 1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _274_
timestamp 1666464484
transform 1 0 19044 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _275_
timestamp 1666464484
transform 1 0 18032 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _276_
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _277_
timestamp 1666464484
transform 1 0 20424 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _278_
timestamp 1666464484
transform -1 0 15180 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1666464484
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1666464484
transform 1 0 8464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _281_
timestamp 1666464484
transform -1 0 14168 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1666464484
transform -1 0 13432 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _283_
timestamp 1666464484
transform 1 0 12696 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _284_
timestamp 1666464484
transform -1 0 15088 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _285_
timestamp 1666464484
transform -1 0 15916 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _286_
timestamp 1666464484
transform -1 0 14996 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1666464484
transform 1 0 8372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _288_
timestamp 1666464484
transform -1 0 12328 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _289_
timestamp 1666464484
transform 1 0 12512 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _290_
timestamp 1666464484
transform -1 0 12788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _291_
timestamp 1666464484
transform 1 0 11684 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _292_
timestamp 1666464484
transform -1 0 10948 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1666464484
transform 1 0 4784 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1666464484
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _295_
timestamp 1666464484
transform 1 0 3956 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1666464484
transform -1 0 3128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _297_
timestamp 1666464484
transform -1 0 4968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _298_
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _299_
timestamp 1666464484
transform 1 0 3956 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _300_
timestamp 1666464484
transform -1 0 4692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1666464484
transform 1 0 3956 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _302_
timestamp 1666464484
transform -1 0 2208 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _303_
timestamp 1666464484
transform -1 0 4048 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _304_
timestamp 1666464484
transform 1 0 2576 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_4  _305_
timestamp 1666464484
transform 1 0 1564 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _306_
timestamp 1666464484
transform 1 0 6532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _307_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14168 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp 1666464484
transform 1 0 10304 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp 1666464484
transform 1 0 7360 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp 1666464484
transform 1 0 7820 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _311_
timestamp 1666464484
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _312_
timestamp 1666464484
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _313_
timestamp 1666464484
transform -1 0 4876 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _314_
timestamp 1666464484
transform -1 0 3036 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _315_
timestamp 1666464484
transform -1 0 3036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _316_
timestamp 1666464484
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _317_
timestamp 1666464484
transform -1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _318_
timestamp 1666464484
transform -1 0 3036 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _319_
timestamp 1666464484
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _320_
timestamp 1666464484
transform -1 0 5336 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _321_
timestamp 1666464484
transform -1 0 3036 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _322_
timestamp 1666464484
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _323_
timestamp 1666464484
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _324_
timestamp 1666464484
transform -1 0 3036 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _325_
timestamp 1666464484
transform -1 0 13156 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1666464484
transform -1 0 11224 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1666464484
transform 1 0 10672 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1666464484
transform -1 0 11224 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1666464484
transform 1 0 9752 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1666464484
transform 1 0 10396 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1666464484
transform 1 0 7176 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1666464484
transform -1 0 21528 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1666464484
transform -1 0 22356 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1666464484
transform -1 0 22356 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _335_
timestamp 1666464484
transform -1 0 21528 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _336_
timestamp 1666464484
transform -1 0 22356 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _337_
timestamp 1666464484
transform 1 0 20884 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _338_
timestamp 1666464484
transform -1 0 21528 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1666464484
transform 1 0 7452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1666464484
transform -1 0 10764 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout31
timestamp 1666464484
transform -1 0 6072 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout32 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 19688 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform -1 0 19412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1666464484
transform -1 0 18032 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform -1 0 20608 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform 1 0 15732 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform -1 0 6072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1666464484
transform -1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform -1 0 5704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1666464484
transform 1 0 4600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1666464484
transform 1 0 7176 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1666464484
transform 1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1666464484
transform -1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1666464484
transform 1 0 5888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1666464484
transform -1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1666464484
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1666464484
transform -1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1666464484
transform -1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1666464484
transform 1 0 3680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1666464484
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1666464484
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1666464484
transform -1 0 22356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1666464484
transform 1 0 22080 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform 1 0 22080 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform 1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform 1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform 1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform 1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform 1 0 22080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform 1 0 22080 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform 1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform 1 0 17940 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform 1 0 18400 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform 1 0 19688 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform -1 0 19688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform -1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform -1 0 14720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform -1 0 11960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform 1 0 6072 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform -1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform -1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform -1 0 6808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform -1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform -1 0 5244 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform -1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform -1 0 3772 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform -1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform -1 0 1840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform -1 0 3312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform 1 0 22080 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform 1 0 22080 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform 1 0 22080 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_78
timestamp 1666464484
transform 1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_79
timestamp 1666464484
transform 1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_80
timestamp 1666464484
transform 1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_81
timestamp 1666464484
transform 1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_82
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_83
timestamp 1666464484
transform 1 0 19780 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_84
timestamp 1666464484
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_85
timestamp 1666464484
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_86
timestamp 1666464484
transform 1 0 19044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_87
timestamp 1666464484
transform -1 0 20332 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_88
timestamp 1666464484
transform -1 0 17756 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_89
timestamp 1666464484
transform -1 0 15364 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_90
timestamp 1666464484
transform 1 0 9108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_91
timestamp 1666464484
transform -1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_92
timestamp 1666464484
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_93
timestamp 1666464484
transform -1 0 4784 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_94
timestamp 1666464484
transform -1 0 6440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_95
timestamp 1666464484
transform -1 0 8096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_96
timestamp 1666464484
transform -1 0 5888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_97
timestamp 1666464484
transform -1 0 5796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_98
timestamp 1666464484
transform -1 0 5520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_99
timestamp 1666464484
transform -1 0 2668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_100
timestamp 1666464484
transform -1 0 3772 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_101
timestamp 1666464484
transform -1 0 5520 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_102
timestamp 1666464484
transform -1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_103
timestamp 1666464484
transform -1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_104
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_105
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_106
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_107
timestamp 1666464484
transform -1 0 1840 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 23200 2864 24000 2984 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 23200 19184 24000 19304 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 23200 20816 24000 20936 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 23200 22448 24000 22568 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 23200 24080 24000 24200 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 23200 25712 24000 25832 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 22742 29200 22798 30000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 20258 29200 20314 30000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 17774 29200 17830 30000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 15290 29200 15346 30000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 12806 29200 12862 30000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 23200 4496 24000 4616 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 10322 29200 10378 30000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 7838 29200 7894 30000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 5354 29200 5410 30000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 2870 29200 2926 30000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 23200 6128 24000 6248 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 23200 7760 24000 7880 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 23200 9392 24000 9512 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 23200 11024 24000 11144 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 23200 12656 24000 12776 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 23200 14288 24000 14408 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 23200 15920 24000 16040 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 23200 17552 24000 17672 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 23200 3952 24000 4072 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 23200 20272 24000 20392 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 23200 21904 24000 22024 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 23200 23536 24000 23656 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 23200 25168 24000 25288 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 23200 26800 24000 26920 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 21086 29200 21142 30000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 18602 29200 18658 30000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 13634 29200 13690 30000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 11150 29200 11206 30000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 23200 5584 24000 5704 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 8666 29200 8722 30000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 6182 29200 6238 30000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 3698 29200 3754 30000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 1214 29200 1270 30000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 23200 7216 24000 7336 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 23200 8848 24000 8968 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 23200 10480 24000 10600 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 23200 12112 24000 12232 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 23200 13744 24000 13864 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 23200 15376 24000 15496 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 23200 17008 24000 17128 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 23200 18640 24000 18760 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 23200 3408 24000 3528 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 23200 19728 24000 19848 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 23200 21360 24000 21480 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 23200 22992 24000 23112 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 23200 24624 24000 24744 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 23200 26256 24000 26376 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 21914 29200 21970 30000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 19430 29200 19486 30000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 16946 29200 17002 30000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 14462 29200 14518 30000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 11978 29200 12034 30000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 23200 5040 24000 5160 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 9494 29200 9550 30000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 7010 29200 7066 30000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 4526 29200 4582 30000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 2042 29200 2098 30000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 23200 6672 24000 6792 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 23200 8304 24000 8424 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 23200 9936 24000 10056 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 23200 11568 24000 11688 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 23200 13200 24000 13320 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 23200 14832 24000 14952 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 23200 16464 24000 16584 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 23200 18096 24000 18216 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 3658 2128 3978 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 9086 2128 9406 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 14514 2128 14834 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 19942 2128 20262 27792 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 6372 2128 6692 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 27792 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 11960 27744 11960 27744 0 vccd1
rlabel via1 12040 27200 12040 27200 0 vssd1
rlabel metal1 14582 20536 14582 20536 0 _000_
rlabel metal1 10396 21862 10396 21862 0 _001_
rlabel metal1 7390 20502 7390 20502 0 _002_
rlabel metal1 7758 18326 7758 18326 0 _003_
rlabel metal2 4462 17374 4462 17374 0 _004_
rlabel metal1 2070 19482 2070 19482 0 _005_
rlabel metal2 6578 15878 6578 15878 0 _006_
rlabel metal2 5934 15912 5934 15912 0 _007_
rlabel metal2 2898 16490 2898 16490 0 _008_
rlabel metal1 1778 17578 1778 17578 0 _009_
rlabel metal1 5382 15096 5382 15096 0 _010_
rlabel via1 2718 25262 2718 25262 0 _011_
rlabel via1 1881 21998 1881 21998 0 _012_
rlabel metal1 4416 21658 4416 21658 0 _013_
rlabel via1 2718 24174 2718 24174 0 _014_
rlabel metal1 2318 23086 2318 23086 0 _015_
rlabel metal1 1877 22712 1877 22712 0 _016_
rlabel via1 2718 24786 2718 24786 0 _017_
rlabel metal1 13028 26962 13028 26962 0 _018_
rlabel metal1 10948 23834 10948 23834 0 _019_
rlabel metal2 10442 25330 10442 25330 0 _020_
rlabel metal1 11822 24922 11822 24922 0 _021_
rlabel metal1 9522 24650 9522 24650 0 _022_
rlabel metal1 10616 25262 10616 25262 0 _023_
rlabel metal2 6946 26962 6946 26962 0 _024_
rlabel metal1 21359 22678 21359 22678 0 _025_
rlabel metal2 22034 24922 22034 24922 0 _026_
rlabel metal1 21624 21998 21624 21998 0 _027_
rlabel metal1 21400 24786 21400 24786 0 _028_
rlabel metal1 21302 25262 21302 25262 0 _029_
rlabel metal1 21104 20910 21104 20910 0 _030_
rlabel metal1 21635 23766 21635 23766 0 _031_
rlabel via2 19550 22933 19550 22933 0 _032_
rlabel metal1 19826 21658 19826 21658 0 _033_
rlabel metal1 18262 23630 18262 23630 0 _034_
rlabel metal1 18998 22406 18998 22406 0 _035_
rlabel metal2 18630 22746 18630 22746 0 _036_
rlabel metal1 20010 22100 20010 22100 0 _037_
rlabel metal1 15962 20366 15962 20366 0 _038_
rlabel metal2 12926 26605 12926 26605 0 _039_
rlabel metal1 12926 26316 12926 26316 0 _040_
rlabel metal1 13340 27098 13340 27098 0 _041_
rlabel metal2 13294 26452 13294 26452 0 _042_
rlabel metal1 13570 26010 13570 26010 0 _043_
rlabel metal2 14582 27302 14582 27302 0 _044_
rlabel metal1 15180 27438 15180 27438 0 _045_
rlabel metal2 13478 26248 13478 26248 0 _046_
rlabel metal2 12742 25840 12742 25840 0 _047_
rlabel metal2 12282 25466 12282 25466 0 _048_
rlabel metal2 12558 25738 12558 25738 0 _049_
rlabel metal1 12696 25262 12696 25262 0 _050_
rlabel via1 10626 22073 10626 22073 0 _051_
rlabel metal1 4830 22066 4830 22066 0 _052_
rlabel metal2 4186 24004 4186 24004 0 _053_
rlabel metal2 2530 23868 2530 23868 0 _054_
rlabel metal2 4186 21165 4186 21165 0 _055_
rlabel metal1 4370 23052 4370 23052 0 _056_
rlabel metal1 4480 23086 4480 23086 0 _057_
rlabel metal2 4646 24106 4646 24106 0 _058_
rlabel metal1 3082 21658 3082 21658 0 _059_
rlabel metal1 3726 26282 3726 26282 0 _060_
rlabel metal2 2162 21284 2162 21284 0 _061_
rlabel metal1 3128 24582 3128 24582 0 _062_
rlabel metal2 2622 22644 2622 22644 0 _063_
rlabel metal1 2116 21590 2116 21590 0 _064_
rlabel metal1 1748 13498 1748 13498 0 _065_
rlabel metal1 3542 12410 3542 12410 0 _066_
rlabel metal1 2300 13498 2300 13498 0 _067_
rlabel metal2 4554 14756 4554 14756 0 _068_
rlabel metal1 1610 18632 1610 18632 0 _069_
rlabel via1 4094 15470 4094 15470 0 _070_
rlabel metal1 4002 15504 4002 15504 0 _071_
rlabel metal1 4692 15674 4692 15674 0 _072_
rlabel metal1 2622 13838 2622 13838 0 _073_
rlabel metal2 3174 15572 3174 15572 0 _074_
rlabel metal1 3772 15130 3772 15130 0 _075_
rlabel metal1 2691 15538 2691 15538 0 _076_
rlabel metal1 2116 18326 2116 18326 0 _077_
rlabel metal1 4968 15130 4968 15130 0 _078_
rlabel metal2 5290 16048 5290 16048 0 _079_
rlabel viali 5282 15402 5282 15402 0 _080_
rlabel via2 2438 19363 2438 19363 0 _081_
rlabel metal1 1794 12852 1794 12852 0 _082_
rlabel metal1 2346 18122 2346 18122 0 _083_
rlabel metal1 2461 14042 2461 14042 0 _084_
rlabel metal1 3726 14314 3726 14314 0 _085_
rlabel metal2 4370 17136 4370 17136 0 _086_
rlabel metal2 6118 16082 6118 16082 0 _087_
rlabel metal1 1978 18190 1978 18190 0 _088_
rlabel metal2 1978 18105 1978 18105 0 _089_
rlabel metal2 3358 18564 3358 18564 0 _090_
rlabel metal2 4002 14314 4002 14314 0 _091_
rlabel metal2 4646 13600 4646 13600 0 _092_
rlabel metal1 1610 12240 1610 12240 0 _093_
rlabel metal2 5566 15436 5566 15436 0 _094_
rlabel metal2 2070 26758 2070 26758 0 _095_
rlabel metal1 3036 21114 3036 21114 0 _096_
rlabel metal1 3120 20774 3120 20774 0 _097_
rlabel metal1 2208 21046 2208 21046 0 _098_
rlabel metal1 3082 22542 3082 22542 0 _099_
rlabel metal1 3450 22406 3450 22406 0 _100_
rlabel metal1 4094 22406 4094 22406 0 _101_
rlabel metal2 2070 25330 2070 25330 0 _102_
rlabel metal1 1794 20570 1794 20570 0 _103_
rlabel metal2 2162 25432 2162 25432 0 _104_
rlabel metal1 4148 21930 4148 21930 0 _105_
rlabel metal1 1978 21352 1978 21352 0 _106_
rlabel via2 2162 21675 2162 21675 0 _107_
rlabel metal2 4646 22678 4646 22678 0 _108_
rlabel metal1 5766 22678 5766 22678 0 _109_
rlabel metal1 5290 22406 5290 22406 0 _110_
rlabel metal1 4692 22134 4692 22134 0 _111_
rlabel metal2 17066 26078 17066 26078 0 _112_
rlabel metal1 13294 25772 13294 25772 0 _113_
rlabel via1 8426 26282 8426 26282 0 _114_
rlabel metal1 9982 26486 9982 26486 0 _115_
rlabel metal2 14306 26401 14306 26401 0 _116_
rlabel metal1 8740 26758 8740 26758 0 _117_
rlabel metal1 9890 24174 9890 24174 0 _118_
rlabel metal1 9706 25262 9706 25262 0 _119_
rlabel metal1 10488 24242 10488 24242 0 _120_
rlabel metal2 12834 25670 12834 25670 0 _121_
rlabel metal1 7636 26350 7636 26350 0 _122_
rlabel metal1 10764 24582 10764 24582 0 _123_
rlabel metal1 9154 24752 9154 24752 0 _124_
rlabel metal2 7406 26656 7406 26656 0 _125_
rlabel metal1 6289 27098 6289 27098 0 _126_
rlabel metal1 7268 25874 7268 25874 0 _127_
rlabel metal1 9844 24650 9844 24650 0 _128_
rlabel metal2 22126 24004 22126 24004 0 _129_
rlabel metal3 21367 20604 21367 20604 0 _130_
rlabel metal1 21122 20570 21122 20570 0 _131_
rlabel metal1 21620 20570 21620 20570 0 _132_
rlabel metal2 19274 24293 19274 24293 0 _133_
rlabel metal1 18975 22746 18975 22746 0 _134_
rlabel metal1 20194 23290 20194 23290 0 _135_
rlabel metal1 21390 25670 21390 25670 0 _136_
rlabel metal1 19872 24378 19872 24378 0 _137_
rlabel metal2 22218 25534 22218 25534 0 _138_
rlabel metal1 19274 21964 19274 21964 0 _139_
rlabel metal1 20562 22202 20562 22202 0 _140_
rlabel metal1 20470 21896 20470 21896 0 _141_
rlabel metal2 17618 24106 17618 24106 0 _142_
rlabel metal1 18408 24038 18408 24038 0 _143_
rlabel metal1 19182 24378 19182 24378 0 _144_
rlabel metal2 22218 23443 22218 23443 0 _145_
rlabel metal1 11454 19346 11454 19346 0 _146_
rlabel metal1 21528 23154 21528 23154 0 _147_
rlabel metal1 19504 23698 19504 23698 0 _148_
rlabel metal2 21298 23290 21298 23290 0 _149_
rlabel metal1 18998 22610 18998 22610 0 _150_
rlabel metal1 22264 20026 22264 20026 0 _151_
rlabel via1 21316 21522 21316 21522 0 _152_
rlabel metal2 22034 19295 22034 19295 0 io_in[10]
rlabel metal2 21390 20349 21390 20349 0 io_in[11]
rlabel metal2 19734 21641 19734 21641 0 io_in[12]
rlabel metal1 17250 24208 17250 24208 0 io_in[13]
rlabel metal1 19320 25874 19320 25874 0 io_in[14]
rlabel metal2 22625 29308 22625 29308 0 io_in[15]
rlabel metal1 20562 27574 20562 27574 0 io_in[16]
rlabel metal1 18170 27438 18170 27438 0 io_in[17]
rlabel metal1 15640 26350 15640 26350 0 io_in[18]
rlabel metal1 13386 26350 13386 26350 0 io_in[19]
rlabel metal2 9982 28203 9982 28203 0 io_in[20]
rlabel metal1 6716 22066 6716 22066 0 io_in[21]
rlabel metal2 5474 25364 5474 25364 0 io_in[22]
rlabel metal1 4830 26282 4830 26282 0 io_in[23]
rlabel metal1 7452 24786 7452 24786 0 io_in[24]
rlabel metal1 6992 25262 6992 25262 0 io_in[25]
rlabel metal3 1602 24820 1602 24820 0 io_in[26]
rlabel metal1 5014 22610 5014 22610 0 io_in[27]
rlabel metal2 3082 20587 3082 20587 0 io_in[28]
rlabel metal1 1564 19822 1564 19822 0 io_in[29]
rlabel metal2 2806 17697 2806 17697 0 io_in[30]
rlabel metal3 1717 14620 1717 14620 0 io_in[31]
rlabel metal1 3726 12818 3726 12818 0 io_in[32]
rlabel metal2 1610 10591 1610 10591 0 io_in[33]
rlabel metal2 1794 8721 1794 8721 0 io_in[34]
rlabel metal2 22126 16031 22126 16031 0 io_in[8]
rlabel via2 22310 17629 22310 17629 0 io_in[9]
rlabel metal3 1188 5780 1188 5780 0 io_out[35]
rlabel metal1 17710 22644 17710 22644 0 mod.clock_counter_a\[0\]
rlabel metal1 17526 22576 17526 22576 0 mod.clock_counter_a\[1\]
rlabel metal1 18446 22644 18446 22644 0 mod.clock_counter_a\[2\]
rlabel metal2 18078 24208 18078 24208 0 mod.clock_counter_a\[3\]
rlabel metal1 20470 21114 20470 21114 0 mod.clock_counter_a\[4\]
rlabel metal2 19090 23358 19090 23358 0 mod.clock_counter_a\[5\]
rlabel metal2 20470 23290 20470 23290 0 mod.clock_counter_a\[6\]
rlabel metal1 14674 26248 14674 26248 0 mod.clock_counter_b\[0\]
rlabel metal1 7866 26928 7866 26928 0 mod.clock_counter_b\[1\]
rlabel metal1 12052 26486 12052 26486 0 mod.clock_counter_b\[2\]
rlabel metal1 8740 25806 8740 25806 0 mod.clock_counter_b\[3\]
rlabel metal1 12834 26384 12834 26384 0 mod.clock_counter_b\[4\]
rlabel metal1 7590 26248 7590 26248 0 mod.clock_counter_b\[5\]
rlabel metal1 11730 27472 11730 27472 0 mod.clock_counter_b\[6\]
rlabel metal2 1610 25874 1610 25874 0 mod.clock_counter_c\[0\]
rlabel metal1 2530 25874 2530 25874 0 mod.clock_counter_c\[1\]
rlabel metal1 1886 20876 1886 20876 0 mod.clock_counter_c\[2\]
rlabel metal1 1702 20910 1702 20910 0 mod.clock_counter_c\[3\]
rlabel metal1 4278 24140 4278 24140 0 mod.clock_counter_c\[4\]
rlabel metal1 3450 21930 3450 21930 0 mod.clock_counter_c\[5\]
rlabel metal2 1610 24140 1610 24140 0 mod.clock_counter_c\[6\]
rlabel metal2 2990 17782 2990 17782 0 mod.clock_counter_d\[0\]
rlabel metal2 3082 18598 3082 18598 0 mod.clock_counter_d\[1\]
rlabel metal1 3404 16218 3404 16218 0 mod.clock_counter_d\[2\]
rlabel metal1 2116 16218 2116 16218 0 mod.clock_counter_d\[3\]
rlabel metal2 2714 13872 2714 13872 0 mod.clock_counter_d\[4\]
rlabel metal2 3082 15521 3082 15521 0 mod.clock_counter_d\[5\]
rlabel metal2 1610 15300 1610 15300 0 mod.clock_counter_d\[6\]
rlabel metal1 9338 15470 9338 15470 0 mod.clock_syn
rlabel metal1 12742 20366 12742 20366 0 mod.div_clock\[0\]
rlabel metal1 13570 19414 13570 19414 0 mod.div_clock\[1\]
rlabel metal2 12558 19788 12558 19788 0 mod.div_clock\[2\]
rlabel metal1 9384 18394 9384 18394 0 mod.div_clock\[3\]
rlabel metal1 12834 19210 12834 19210 0 net1
rlabel metal2 13386 25738 13386 25738 0 net10
rlabel via2 3542 18037 3542 18037 0 net100
rlabel metal2 4186 16507 4186 16507 0 net101
rlabel metal2 3910 14161 3910 14161 0 net102
rlabel metal2 2254 11815 2254 11815 0 net103
rlabel metal3 1142 9860 1142 9860 0 net104
rlabel metal3 1142 7820 1142 7820 0 net105
rlabel metal3 1142 3740 1142 3740 0 net106
rlabel metal3 1142 1700 1142 1700 0 net107
rlabel metal1 8464 25262 8464 25262 0 net11
rlabel metal1 8418 24786 8418 24786 0 net12
rlabel metal2 7774 25874 7774 25874 0 net13
rlabel metal1 4646 26452 4646 26452 0 net14
rlabel metal1 5014 24786 5014 24786 0 net15
rlabel metal1 6578 25466 6578 25466 0 net16
rlabel metal2 2438 26826 2438 26826 0 net17
rlabel metal2 5934 23494 5934 23494 0 net18
rlabel metal1 4048 20570 4048 20570 0 net19
rlabel metal1 21022 20026 21022 20026 0 net2
rlabel metal2 3450 18428 3450 18428 0 net20
rlabel metal1 2070 18802 2070 18802 0 net21
rlabel metal1 4324 13498 4324 13498 0 net22
rlabel metal1 1794 11764 1794 11764 0 net23
rlabel metal1 2300 10778 2300 10778 0 net24
rlabel metal1 1564 9146 1564 9146 0 net25
rlabel metal1 22218 22610 22218 22610 0 net26
rlabel metal1 22172 17850 22172 17850 0 net27
rlabel metal1 4692 6290 4692 6290 0 net28
rlabel metal1 16008 26826 16008 26826 0 net29
rlabel metal2 19642 20332 19642 20332 0 net3
rlabel metal1 1610 16694 1610 16694 0 net30
rlabel metal1 12558 27608 12558 27608 0 net31
rlabel metal1 22310 21964 22310 21964 0 net32
rlabel via2 22310 3995 22310 3995 0 net33
rlabel via2 22310 5661 22310 5661 0 net34
rlabel via2 22310 7259 22310 7259 0 net35
rlabel via2 22310 8925 22310 8925 0 net36
rlabel via2 22310 10523 22310 10523 0 net37
rlabel via2 22310 12189 22310 12189 0 net38
rlabel via2 22310 13821 22310 13821 0 net39
rlabel metal2 17434 24582 17434 24582 0 net4
rlabel via2 22310 15453 22310 15453 0 net40
rlabel via2 22310 17051 22310 17051 0 net41
rlabel via2 22310 18717 22310 18717 0 net42
rlabel metal2 22034 20825 22034 20825 0 net43
rlabel metal1 20562 20434 20562 20434 0 net44
rlabel metal2 19826 24123 19826 24123 0 net45
rlabel metal2 20654 25789 20654 25789 0 net46
rlabel via2 20562 26877 20562 26877 0 net47
rlabel metal1 20516 26826 20516 26826 0 net48
rlabel metal1 19044 27438 19044 27438 0 net49
rlabel metal2 22126 26588 22126 26588 0 net5
rlabel metal1 16744 26962 16744 26962 0 net50
rlabel metal1 14214 25806 14214 25806 0 net51
rlabel metal1 11454 24378 11454 24378 0 net52
rlabel metal1 7498 26418 7498 26418 0 net53
rlabel metal1 6394 25874 6394 25874 0 net54
rlabel metal1 3680 26962 3680 26962 0 net55
rlabel metal2 1242 27329 1242 27329 0 net56
rlabel metal1 7268 24310 7268 24310 0 net57
rlabel metal2 3450 25619 3450 25619 0 net58
rlabel metal2 2898 25109 2898 25109 0 net59
rlabel metal1 19550 26384 19550 26384 0 net6
rlabel via2 3174 21437 3174 21437 0 net60
rlabel metal3 1464 19380 1464 19380 0 net61
rlabel metal3 1142 17340 1142 17340 0 net62
rlabel metal2 3082 14059 3082 14059 0 net63
rlabel metal1 2530 12410 2530 12410 0 net64
rlabel metal3 1786 11220 1786 11220 0 net65
rlabel metal3 1142 9180 1142 9180 0 net66
rlabel metal3 1142 7140 1142 7140 0 net67
rlabel metal3 1142 5100 1142 5100 0 net68
rlabel metal3 1142 3060 1142 3060 0 net69
rlabel metal2 20562 27268 20562 27268 0 net7
rlabel metal3 1050 1020 1050 1020 0 net70
rlabel via2 22310 3485 22310 3485 0 net71
rlabel via2 22310 5083 22310 5083 0 net72
rlabel via2 22310 6749 22310 6749 0 net73
rlabel via2 22310 8347 22310 8347 0 net74
rlabel via2 22310 10013 22310 10013 0 net75
rlabel via2 22310 11611 22310 11611 0 net76
rlabel via2 22310 13277 22310 13277 0 net77
rlabel via2 22310 14875 22310 14875 0 net78
rlabel metal2 22034 16575 22034 16575 0 net79
rlabel metal1 16606 27030 16606 27030 0 net8
rlabel via2 22310 18139 22310 18139 0 net80
rlabel metal2 22310 20009 22310 20009 0 net81
rlabel via2 19458 21437 19458 21437 0 net82
rlabel metal1 20194 20434 20194 20434 0 net83
rlabel metal2 21482 25721 21482 25721 0 net84
rlabel via2 19458 26333 19458 26333 0 net85
rlabel metal1 19274 26996 19274 26996 0 net86
rlabel metal1 19780 27574 19780 27574 0 net87
rlabel metal1 17250 27574 17250 27574 0 net88
rlabel metal1 14766 26486 14766 26486 0 net89
rlabel metal2 15778 26078 15778 26078 0 net9
rlabel metal1 10672 27642 10672 27642 0 net90
rlabel metal2 9614 26843 9614 26843 0 net91
rlabel metal1 5796 27574 5796 27574 0 net92
rlabel metal2 4554 28128 4554 28128 0 net93
rlabel metal2 2215 29308 2215 29308 0 net94
rlabel metal1 7728 24786 7728 24786 0 net95
rlabel metal1 4876 25806 4876 25806 0 net96
rlabel metal2 4094 24412 4094 24412 0 net97
rlabel metal3 1717 22100 1717 22100 0 net98
rlabel metal3 1556 20060 1556 20060 0 net99
<< properties >>
string FIXED_BBOX 0 0 24000 30000
<< end >>
