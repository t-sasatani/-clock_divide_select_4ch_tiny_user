magic
tech sky130A
magscale 1 2
timestamp 1672331279
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 2128 58880 57712
<< metal2 >>
rect 1214 59200 1270 60000
rect 3422 59200 3478 60000
rect 5630 59200 5686 60000
rect 7838 59200 7894 60000
rect 10046 59200 10102 60000
rect 12254 59200 12310 60000
rect 14462 59200 14518 60000
rect 16670 59200 16726 60000
rect 18878 59200 18934 60000
rect 21086 59200 21142 60000
rect 23294 59200 23350 60000
rect 25502 59200 25558 60000
rect 27710 59200 27766 60000
rect 29918 59200 29974 60000
rect 32126 59200 32182 60000
rect 34334 59200 34390 60000
rect 36542 59200 36598 60000
rect 38750 59200 38806 60000
rect 40958 59200 41014 60000
rect 43166 59200 43222 60000
rect 45374 59200 45430 60000
rect 47582 59200 47638 60000
rect 49790 59200 49846 60000
rect 51998 59200 52054 60000
rect 54206 59200 54262 60000
rect 56414 59200 56470 60000
rect 58622 59200 58678 60000
<< obsm2 >>
rect 1326 59144 3366 59200
rect 3534 59144 5574 59200
rect 5742 59144 7782 59200
rect 7950 59144 9990 59200
rect 10158 59144 12198 59200
rect 12366 59144 14406 59200
rect 14574 59144 16614 59200
rect 16782 59144 18822 59200
rect 18990 59144 21030 59200
rect 21198 59144 23238 59200
rect 23406 59144 25446 59200
rect 25614 59144 27654 59200
rect 27822 59144 29862 59200
rect 30030 59144 32070 59200
rect 32238 59144 34278 59200
rect 34446 59144 36486 59200
rect 36654 59144 38694 59200
rect 38862 59144 40902 59200
rect 41070 59144 43110 59200
rect 43278 59144 45318 59200
rect 45486 59144 47526 59200
rect 47694 59144 49734 59200
rect 49902 59144 51942 59200
rect 52110 59144 54150 59200
rect 54318 59144 56358 59200
rect 56526 59144 58402 59200
rect 1216 2071 58402 59144
<< metal3 >>
rect 0 57808 800 57928
rect 59200 56856 60000 56976
rect 0 56448 800 56568
rect 59200 55632 60000 55752
rect 0 55088 800 55208
rect 59200 54408 60000 54528
rect 0 53728 800 53848
rect 59200 53184 60000 53304
rect 0 52368 800 52488
rect 59200 51960 60000 52080
rect 0 51008 800 51128
rect 59200 50736 60000 50856
rect 0 49648 800 49768
rect 59200 49512 60000 49632
rect 0 48288 800 48408
rect 59200 48288 60000 48408
rect 0 46928 800 47048
rect 59200 47064 60000 47184
rect 59200 45840 60000 45960
rect 0 45568 800 45688
rect 59200 44616 60000 44736
rect 0 44208 800 44328
rect 59200 43392 60000 43512
rect 0 42848 800 42968
rect 59200 42168 60000 42288
rect 0 41488 800 41608
rect 59200 40944 60000 41064
rect 0 40128 800 40248
rect 59200 39720 60000 39840
rect 0 38768 800 38888
rect 59200 38496 60000 38616
rect 0 37408 800 37528
rect 59200 37272 60000 37392
rect 0 36048 800 36168
rect 59200 36048 60000 36168
rect 0 34688 800 34808
rect 59200 34824 60000 34944
rect 59200 33600 60000 33720
rect 0 33328 800 33448
rect 59200 32376 60000 32496
rect 0 31968 800 32088
rect 59200 31152 60000 31272
rect 0 30608 800 30728
rect 59200 29928 60000 30048
rect 0 29248 800 29368
rect 59200 28704 60000 28824
rect 0 27888 800 28008
rect 59200 27480 60000 27600
rect 0 26528 800 26648
rect 59200 26256 60000 26376
rect 0 25168 800 25288
rect 59200 25032 60000 25152
rect 0 23808 800 23928
rect 59200 23808 60000 23928
rect 0 22448 800 22568
rect 59200 22584 60000 22704
rect 59200 21360 60000 21480
rect 0 21088 800 21208
rect 59200 20136 60000 20256
rect 0 19728 800 19848
rect 59200 18912 60000 19032
rect 0 18368 800 18488
rect 59200 17688 60000 17808
rect 0 17008 800 17128
rect 59200 16464 60000 16584
rect 0 15648 800 15768
rect 59200 15240 60000 15360
rect 0 14288 800 14408
rect 59200 14016 60000 14136
rect 0 12928 800 13048
rect 59200 12792 60000 12912
rect 0 11568 800 11688
rect 59200 11568 60000 11688
rect 0 10208 800 10328
rect 59200 10344 60000 10464
rect 59200 9120 60000 9240
rect 0 8848 800 8968
rect 59200 7896 60000 8016
rect 0 7488 800 7608
rect 59200 6672 60000 6792
rect 0 6128 800 6248
rect 59200 5448 60000 5568
rect 0 4768 800 4888
rect 59200 4224 60000 4344
rect 0 3408 800 3528
rect 59200 3000 60000 3120
rect 0 2048 800 2168
<< obsm3 >>
rect 800 57056 59200 57697
rect 800 56776 59120 57056
rect 800 56648 59200 56776
rect 880 56368 59200 56648
rect 800 55832 59200 56368
rect 800 55552 59120 55832
rect 800 55288 59200 55552
rect 880 55008 59200 55288
rect 800 54608 59200 55008
rect 800 54328 59120 54608
rect 800 53928 59200 54328
rect 880 53648 59200 53928
rect 800 53384 59200 53648
rect 800 53104 59120 53384
rect 800 52568 59200 53104
rect 880 52288 59200 52568
rect 800 52160 59200 52288
rect 800 51880 59120 52160
rect 800 51208 59200 51880
rect 880 50936 59200 51208
rect 880 50928 59120 50936
rect 800 50656 59120 50928
rect 800 49848 59200 50656
rect 880 49712 59200 49848
rect 880 49568 59120 49712
rect 800 49432 59120 49568
rect 800 48488 59200 49432
rect 880 48208 59120 48488
rect 800 47264 59200 48208
rect 800 47128 59120 47264
rect 880 46984 59120 47128
rect 880 46848 59200 46984
rect 800 46040 59200 46848
rect 800 45768 59120 46040
rect 880 45760 59120 45768
rect 880 45488 59200 45760
rect 800 44816 59200 45488
rect 800 44536 59120 44816
rect 800 44408 59200 44536
rect 880 44128 59200 44408
rect 800 43592 59200 44128
rect 800 43312 59120 43592
rect 800 43048 59200 43312
rect 880 42768 59200 43048
rect 800 42368 59200 42768
rect 800 42088 59120 42368
rect 800 41688 59200 42088
rect 880 41408 59200 41688
rect 800 41144 59200 41408
rect 800 40864 59120 41144
rect 800 40328 59200 40864
rect 880 40048 59200 40328
rect 800 39920 59200 40048
rect 800 39640 59120 39920
rect 800 38968 59200 39640
rect 880 38696 59200 38968
rect 880 38688 59120 38696
rect 800 38416 59120 38688
rect 800 37608 59200 38416
rect 880 37472 59200 37608
rect 880 37328 59120 37472
rect 800 37192 59120 37328
rect 800 36248 59200 37192
rect 880 35968 59120 36248
rect 800 35024 59200 35968
rect 800 34888 59120 35024
rect 880 34744 59120 34888
rect 880 34608 59200 34744
rect 800 33800 59200 34608
rect 800 33528 59120 33800
rect 880 33520 59120 33528
rect 880 33248 59200 33520
rect 800 32576 59200 33248
rect 800 32296 59120 32576
rect 800 32168 59200 32296
rect 880 31888 59200 32168
rect 800 31352 59200 31888
rect 800 31072 59120 31352
rect 800 30808 59200 31072
rect 880 30528 59200 30808
rect 800 30128 59200 30528
rect 800 29848 59120 30128
rect 800 29448 59200 29848
rect 880 29168 59200 29448
rect 800 28904 59200 29168
rect 800 28624 59120 28904
rect 800 28088 59200 28624
rect 880 27808 59200 28088
rect 800 27680 59200 27808
rect 800 27400 59120 27680
rect 800 26728 59200 27400
rect 880 26456 59200 26728
rect 880 26448 59120 26456
rect 800 26176 59120 26448
rect 800 25368 59200 26176
rect 880 25232 59200 25368
rect 880 25088 59120 25232
rect 800 24952 59120 25088
rect 800 24008 59200 24952
rect 880 23728 59120 24008
rect 800 22784 59200 23728
rect 800 22648 59120 22784
rect 880 22504 59120 22648
rect 880 22368 59200 22504
rect 800 21560 59200 22368
rect 800 21288 59120 21560
rect 880 21280 59120 21288
rect 880 21008 59200 21280
rect 800 20336 59200 21008
rect 800 20056 59120 20336
rect 800 19928 59200 20056
rect 880 19648 59200 19928
rect 800 19112 59200 19648
rect 800 18832 59120 19112
rect 800 18568 59200 18832
rect 880 18288 59200 18568
rect 800 17888 59200 18288
rect 800 17608 59120 17888
rect 800 17208 59200 17608
rect 880 16928 59200 17208
rect 800 16664 59200 16928
rect 800 16384 59120 16664
rect 800 15848 59200 16384
rect 880 15568 59200 15848
rect 800 15440 59200 15568
rect 800 15160 59120 15440
rect 800 14488 59200 15160
rect 880 14216 59200 14488
rect 880 14208 59120 14216
rect 800 13936 59120 14208
rect 800 13128 59200 13936
rect 880 12992 59200 13128
rect 880 12848 59120 12992
rect 800 12712 59120 12848
rect 800 11768 59200 12712
rect 880 11488 59120 11768
rect 800 10544 59200 11488
rect 800 10408 59120 10544
rect 880 10264 59120 10408
rect 880 10128 59200 10264
rect 800 9320 59200 10128
rect 800 9048 59120 9320
rect 880 9040 59120 9048
rect 880 8768 59200 9040
rect 800 8096 59200 8768
rect 800 7816 59120 8096
rect 800 7688 59200 7816
rect 880 7408 59200 7688
rect 800 6872 59200 7408
rect 800 6592 59120 6872
rect 800 6328 59200 6592
rect 880 6048 59200 6328
rect 800 5648 59200 6048
rect 800 5368 59120 5648
rect 800 4968 59200 5368
rect 880 4688 59200 4968
rect 800 4424 59200 4688
rect 800 4144 59120 4424
rect 800 3608 59200 4144
rect 880 3328 59200 3608
rect 800 3200 59200 3328
rect 800 2920 59120 3200
rect 800 2248 59200 2920
rect 880 2075 59200 2248
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal3 s 59200 3000 60000 3120 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 59200 39720 60000 39840 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 59200 43392 60000 43512 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 59200 47064 60000 47184 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 59200 50736 60000 50856 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 59200 54408 60000 54528 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 58622 59200 58678 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 51998 59200 52054 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 45374 59200 45430 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 38750 59200 38806 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 32126 59200 32182 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 59200 6672 60000 6792 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 25502 59200 25558 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 18878 59200 18934 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 12254 59200 12310 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 5630 59200 5686 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 59200 10344 60000 10464 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 59200 14016 60000 14136 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59200 17688 60000 17808 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 59200 21360 60000 21480 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 59200 25032 60000 25152 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 59200 28704 60000 28824 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 59200 32376 60000 32496 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 59200 36048 60000 36168 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 59200 5448 60000 5568 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 59200 45840 60000 45960 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 59200 49512 60000 49632 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 59200 53184 60000 53304 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 59200 56856 60000 56976 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 54206 59200 54262 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 47582 59200 47638 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 40958 59200 41014 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 34334 59200 34390 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 27710 59200 27766 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 59200 9120 60000 9240 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 21086 59200 21142 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 14462 59200 14518 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 7838 59200 7894 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 1214 59200 1270 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 59200 16464 60000 16584 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 59200 20136 60000 20256 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 59200 23808 60000 23928 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 59200 27480 60000 27600 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 59200 31152 60000 31272 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 59200 34824 60000 34944 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 59200 38496 60000 38616 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 59200 4224 60000 4344 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 59200 40944 60000 41064 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 59200 44616 60000 44736 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 59200 48288 60000 48408 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 59200 51960 60000 52080 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 59200 55632 60000 55752 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 56414 59200 56470 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 49790 59200 49846 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 43166 59200 43222 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 36542 59200 36598 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 29918 59200 29974 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 23294 59200 23350 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 16670 59200 16726 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 10046 59200 10102 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 3422 59200 3478 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 59200 11568 60000 11688 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 59200 15240 60000 15360 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 59200 18912 60000 19032 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 59200 26256 60000 26376 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 59200 29928 60000 30048 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 59200 33600 60000 33720 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 59200 37272 60000 37392 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 968468
string GDS_FILE /home/runner/work/clock_divide_select_4ch_tiny_user/clock_divide_select_4ch_tiny_user/openlane/tiny_user_project/runs/22_12_29_16_26/results/signoff/tiny_user_project.magic.gds
string GDS_START 23768
<< end >>

