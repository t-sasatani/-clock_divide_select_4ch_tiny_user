// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire net34;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net35;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net36;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net72;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net73;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net74;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire \mod.clock_counter_a[0] ;
 wire \mod.clock_counter_a[1] ;
 wire \mod.clock_counter_a[2] ;
 wire \mod.clock_counter_a[3] ;
 wire \mod.clock_counter_a[4] ;
 wire \mod.clock_counter_a[5] ;
 wire \mod.clock_counter_a[6] ;
 wire \mod.clock_counter_b[0] ;
 wire \mod.clock_counter_b[1] ;
 wire \mod.clock_counter_b[2] ;
 wire \mod.clock_counter_b[3] ;
 wire \mod.clock_counter_b[4] ;
 wire \mod.clock_counter_b[5] ;
 wire \mod.clock_counter_b[6] ;
 wire \mod.clock_counter_c[0] ;
 wire \mod.clock_counter_c[1] ;
 wire \mod.clock_counter_c[2] ;
 wire \mod.clock_counter_c[3] ;
 wire \mod.clock_counter_c[4] ;
 wire \mod.clock_counter_c[5] ;
 wire \mod.clock_counter_c[6] ;
 wire \mod.clock_counter_d[0] ;
 wire \mod.clock_counter_d[1] ;
 wire \mod.clock_counter_d[2] ;
 wire \mod.clock_counter_d[3] ;
 wire \mod.clock_counter_d[4] ;
 wire \mod.clock_counter_d[5] ;
 wire \mod.clock_counter_d[6] ;
 wire \mod.clock_syn ;
 wire \mod.div_clock[0] ;
 wire \mod.div_clock[1] ;
 wire \mod.div_clock[2] ;
 wire \mod.div_clock[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;

 sky130_fd_sc_hd__inv_2 _153_ (.A(net25),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _154_ (.A(net24),
    .Y(_066_));
 sky130_fd_sc_hd__o22a_1 _155_ (.A1(\mod.clock_counter_d[5] ),
    .A2(_065_),
    .B1(_066_),
    .B2(\mod.clock_counter_d[4] ),
    .X(_067_));
 sky130_fd_sc_hd__inv_2 _156_ (.A(net22),
    .Y(_068_));
 sky130_fd_sc_hd__or2b_1 _157_ (.A(\mod.clock_counter_d[1] ),
    .B_N(net21),
    .X(_069_));
 sky130_fd_sc_hd__and2b_1 _158_ (.A_N(net20),
    .B(\mod.clock_counter_d[0] ),
    .X(_070_));
 sky130_fd_sc_hd__and2b_1 _159_ (.A_N(net21),
    .B(\mod.clock_counter_d[1] ),
    .X(_071_));
 sky130_fd_sc_hd__a221o_1 _160_ (.A1(\mod.clock_counter_d[2] ),
    .A2(_068_),
    .B1(_069_),
    .B2(_070_),
    .C1(_071_),
    .X(_072_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(net23),
    .Y(_073_));
 sky130_fd_sc_hd__o22a_1 _162_ (.A1(\mod.clock_counter_d[3] ),
    .A2(_073_),
    .B1(_068_),
    .B2(\mod.clock_counter_d[2] ),
    .X(_074_));
 sky130_fd_sc_hd__a22o_1 _163_ (.A1(\mod.clock_counter_d[4] ),
    .A2(_066_),
    .B1(_073_),
    .B2(\mod.clock_counter_d[3] ),
    .X(_075_));
 sky130_fd_sc_hd__a21o_1 _164_ (.A1(_072_),
    .A2(_074_),
    .B1(_075_),
    .X(_076_));
 sky130_fd_sc_hd__a221oi_4 _165_ (.A1(\mod.clock_counter_d[5] ),
    .A2(_065_),
    .B1(_067_),
    .B2(_076_),
    .C1(\mod.clock_counter_d[6] ),
    .Y(_077_));
 sky130_fd_sc_hd__xnor2_1 _166_ (.A(\mod.div_clock[3] ),
    .B(_077_),
    .Y(_003_));
 sky130_fd_sc_hd__and2b_1 _167_ (.A_N(\mod.clock_counter_d[0] ),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_1 _168_ (.A(_078_),
    .X(_004_));
 sky130_fd_sc_hd__or2_1 _169_ (.A(\mod.clock_counter_d[0] ),
    .B(\mod.clock_counter_d[1] ),
    .X(_079_));
 sky130_fd_sc_hd__nand2_1 _170_ (.A(\mod.clock_counter_d[0] ),
    .B(\mod.clock_counter_d[1] ),
    .Y(_080_));
 sky130_fd_sc_hd__and3_1 _171_ (.A(_077_),
    .B(_079_),
    .C(_080_),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(_081_),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _173_ (.A(\mod.clock_counter_d[0] ),
    .B(\mod.clock_counter_d[1] ),
    .C(\mod.clock_counter_d[2] ),
    .X(_082_));
 sky130_fd_sc_hd__a21o_1 _174_ (.A1(\mod.clock_counter_d[0] ),
    .A2(\mod.clock_counter_d[1] ),
    .B1(\mod.clock_counter_d[2] ),
    .X(_083_));
 sky130_fd_sc_hd__and3b_1 _175_ (.A_N(_082_),
    .B(_083_),
    .C(_077_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_1 _176_ (.A(_084_),
    .X(_006_));
 sky130_fd_sc_hd__and2_1 _177_ (.A(\mod.clock_counter_d[3] ),
    .B(_082_),
    .X(_085_));
 sky130_fd_sc_hd__or2_1 _178_ (.A(\mod.clock_counter_d[3] ),
    .B(_082_),
    .X(_086_));
 sky130_fd_sc_hd__and3b_1 _179_ (.A_N(_085_),
    .B(_086_),
    .C(_077_),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_1 _180_ (.A(_087_),
    .X(_007_));
 sky130_fd_sc_hd__and3_1 _181_ (.A(\mod.clock_counter_d[3] ),
    .B(\mod.clock_counter_d[4] ),
    .C(_082_),
    .X(_088_));
 sky130_fd_sc_hd__or2_1 _182_ (.A(\mod.clock_counter_d[4] ),
    .B(_085_),
    .X(_089_));
 sky130_fd_sc_hd__and3b_1 _183_ (.A_N(_088_),
    .B(_089_),
    .C(_077_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(_090_),
    .X(_008_));
 sky130_fd_sc_hd__or2_1 _185_ (.A(\mod.clock_counter_d[5] ),
    .B(_088_),
    .X(_091_));
 sky130_fd_sc_hd__nand2_1 _186_ (.A(\mod.clock_counter_d[5] ),
    .B(_088_),
    .Y(_092_));
 sky130_fd_sc_hd__and3_1 _187_ (.A(_077_),
    .B(_091_),
    .C(_092_),
    .X(_093_));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(_093_),
    .X(_009_));
 sky130_fd_sc_hd__and3_1 _189_ (.A(\mod.clock_counter_d[5] ),
    .B(_077_),
    .C(_088_),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(_094_),
    .X(_010_));
 sky130_fd_sc_hd__and2b_1 _191_ (.A_N(\mod.clock_counter_c[0] ),
    .B(_064_),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(_095_),
    .X(_011_));
 sky130_fd_sc_hd__or2_1 _193_ (.A(\mod.clock_counter_c[0] ),
    .B(\mod.clock_counter_c[1] ),
    .X(_096_));
 sky130_fd_sc_hd__nand2_1 _194_ (.A(\mod.clock_counter_c[0] ),
    .B(\mod.clock_counter_c[1] ),
    .Y(_097_));
 sky130_fd_sc_hd__and3_1 _195_ (.A(_064_),
    .B(_096_),
    .C(_097_),
    .X(_098_));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(_098_),
    .X(_012_));
 sky130_fd_sc_hd__and3_1 _197_ (.A(\mod.clock_counter_c[0] ),
    .B(\mod.clock_counter_c[1] ),
    .C(\mod.clock_counter_c[2] ),
    .X(_099_));
 sky130_fd_sc_hd__a21o_1 _198_ (.A1(\mod.clock_counter_c[0] ),
    .A2(\mod.clock_counter_c[1] ),
    .B1(\mod.clock_counter_c[2] ),
    .X(_100_));
 sky130_fd_sc_hd__and3b_1 _199_ (.A_N(_099_),
    .B(_100_),
    .C(_064_),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(_101_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _201_ (.A(\mod.clock_counter_c[3] ),
    .B(_099_),
    .X(_102_));
 sky130_fd_sc_hd__or2_1 _202_ (.A(\mod.clock_counter_c[3] ),
    .B(_099_),
    .X(_103_));
 sky130_fd_sc_hd__and3b_1 _203_ (.A_N(_102_),
    .B(_103_),
    .C(_064_),
    .X(_104_));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(_104_),
    .X(_014_));
 sky130_fd_sc_hd__and3_1 _205_ (.A(\mod.clock_counter_c[3] ),
    .B(\mod.clock_counter_c[4] ),
    .C(_099_),
    .X(_105_));
 sky130_fd_sc_hd__or2_1 _206_ (.A(\mod.clock_counter_c[4] ),
    .B(_102_),
    .X(_106_));
 sky130_fd_sc_hd__and3b_1 _207_ (.A_N(_105_),
    .B(_106_),
    .C(_064_),
    .X(_107_));
 sky130_fd_sc_hd__clkbuf_1 _208_ (.A(_107_),
    .X(_015_));
 sky130_fd_sc_hd__or2_1 _209_ (.A(\mod.clock_counter_c[5] ),
    .B(_105_),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(\mod.clock_counter_c[5] ),
    .B(_105_),
    .Y(_109_));
 sky130_fd_sc_hd__and3_1 _211_ (.A(_064_),
    .B(_108_),
    .C(_109_),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_1 _212_ (.A(_110_),
    .X(_016_));
 sky130_fd_sc_hd__and3_1 _213_ (.A(\mod.clock_counter_c[5] ),
    .B(_064_),
    .C(_105_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _214_ (.A(_111_),
    .X(_017_));
 sky130_fd_sc_hd__and2b_1 _215_ (.A_N(\mod.clock_counter_b[0] ),
    .B(_051_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _216_ (.A(_112_),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _217_ (.A(\mod.clock_counter_b[0] ),
    .B(\mod.clock_counter_b[1] ),
    .X(_113_));
 sky130_fd_sc_hd__nand2_1 _218_ (.A(\mod.clock_counter_b[0] ),
    .B(\mod.clock_counter_b[1] ),
    .Y(_114_));
 sky130_fd_sc_hd__and3_1 _219_ (.A(_051_),
    .B(_113_),
    .C(_114_),
    .X(_115_));
 sky130_fd_sc_hd__clkbuf_1 _220_ (.A(_115_),
    .X(_019_));
 sky130_fd_sc_hd__and3_1 _221_ (.A(\mod.clock_counter_b[0] ),
    .B(\mod.clock_counter_b[1] ),
    .C(\mod.clock_counter_b[2] ),
    .X(_116_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(\mod.clock_counter_b[0] ),
    .A2(\mod.clock_counter_b[1] ),
    .B1(\mod.clock_counter_b[2] ),
    .X(_117_));
 sky130_fd_sc_hd__and3b_1 _223_ (.A_N(_116_),
    .B(_117_),
    .C(_051_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_1 _224_ (.A(_118_),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _225_ (.A(\mod.clock_counter_b[3] ),
    .B(_116_),
    .X(_119_));
 sky130_fd_sc_hd__or2_1 _226_ (.A(\mod.clock_counter_b[3] ),
    .B(_116_),
    .X(_120_));
 sky130_fd_sc_hd__and3b_1 _227_ (.A_N(_119_),
    .B(_120_),
    .C(_051_),
    .X(_121_));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(_121_),
    .X(_021_));
 sky130_fd_sc_hd__and3_1 _229_ (.A(\mod.clock_counter_b[3] ),
    .B(\mod.clock_counter_b[4] ),
    .C(_116_),
    .X(_122_));
 sky130_fd_sc_hd__or2_1 _230_ (.A(\mod.clock_counter_b[4] ),
    .B(_119_),
    .X(_123_));
 sky130_fd_sc_hd__and3b_1 _231_ (.A_N(_122_),
    .B(_123_),
    .C(_051_),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _232_ (.A(_124_),
    .X(_022_));
 sky130_fd_sc_hd__or2_1 _233_ (.A(\mod.clock_counter_b[5] ),
    .B(_122_),
    .X(_125_));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(\mod.clock_counter_b[5] ),
    .B(_122_),
    .Y(_126_));
 sky130_fd_sc_hd__and3_1 _235_ (.A(_051_),
    .B(_125_),
    .C(_126_),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(_127_),
    .X(_023_));
 sky130_fd_sc_hd__and3_1 _237_ (.A(\mod.clock_counter_b[5] ),
    .B(_051_),
    .C(_122_),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _238_ (.A(_128_),
    .X(_024_));
 sky130_fd_sc_hd__and2b_1 _239_ (.A_N(\mod.clock_counter_a[0] ),
    .B(_038_),
    .X(_129_));
 sky130_fd_sc_hd__clkbuf_1 _240_ (.A(_129_),
    .X(_025_));
 sky130_fd_sc_hd__or2_1 _241_ (.A(\mod.clock_counter_a[0] ),
    .B(\mod.clock_counter_a[1] ),
    .X(_130_));
 sky130_fd_sc_hd__nand2_1 _242_ (.A(\mod.clock_counter_a[0] ),
    .B(\mod.clock_counter_a[1] ),
    .Y(_131_));
 sky130_fd_sc_hd__and3_1 _243_ (.A(_038_),
    .B(_130_),
    .C(_131_),
    .X(_132_));
 sky130_fd_sc_hd__clkbuf_1 _244_ (.A(_132_),
    .X(_026_));
 sky130_fd_sc_hd__and3_1 _245_ (.A(\mod.clock_counter_a[0] ),
    .B(\mod.clock_counter_a[1] ),
    .C(\mod.clock_counter_a[2] ),
    .X(_133_));
 sky130_fd_sc_hd__a21o_1 _246_ (.A1(\mod.clock_counter_a[0] ),
    .A2(\mod.clock_counter_a[1] ),
    .B1(\mod.clock_counter_a[2] ),
    .X(_134_));
 sky130_fd_sc_hd__and3b_1 _247_ (.A_N(_133_),
    .B(_134_),
    .C(_038_),
    .X(_135_));
 sky130_fd_sc_hd__clkbuf_1 _248_ (.A(_135_),
    .X(_027_));
 sky130_fd_sc_hd__and2_1 _249_ (.A(\mod.clock_counter_a[3] ),
    .B(_133_),
    .X(_136_));
 sky130_fd_sc_hd__or2_1 _250_ (.A(\mod.clock_counter_a[3] ),
    .B(_133_),
    .X(_137_));
 sky130_fd_sc_hd__and3b_1 _251_ (.A_N(_136_),
    .B(_137_),
    .C(_038_),
    .X(_138_));
 sky130_fd_sc_hd__clkbuf_1 _252_ (.A(_138_),
    .X(_028_));
 sky130_fd_sc_hd__and3_1 _253_ (.A(\mod.clock_counter_a[3] ),
    .B(\mod.clock_counter_a[4] ),
    .C(_133_),
    .X(_139_));
 sky130_fd_sc_hd__or2_1 _254_ (.A(\mod.clock_counter_a[4] ),
    .B(_136_),
    .X(_140_));
 sky130_fd_sc_hd__and3b_1 _255_ (.A_N(_139_),
    .B(_140_),
    .C(_038_),
    .X(_141_));
 sky130_fd_sc_hd__clkbuf_1 _256_ (.A(_141_),
    .X(_029_));
 sky130_fd_sc_hd__or2_1 _257_ (.A(\mod.clock_counter_a[5] ),
    .B(_139_),
    .X(_142_));
 sky130_fd_sc_hd__nand2_1 _258_ (.A(\mod.clock_counter_a[5] ),
    .B(_139_),
    .Y(_143_));
 sky130_fd_sc_hd__and3_1 _259_ (.A(_038_),
    .B(_142_),
    .C(_143_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_144_),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _261_ (.A(\mod.clock_counter_a[5] ),
    .B(_038_),
    .C(_139_),
    .X(_145_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_145_),
    .X(_031_));
 sky130_fd_sc_hd__mux4_1 _263_ (.A0(\mod.div_clock[0] ),
    .A1(\mod.div_clock[1] ),
    .A2(\mod.div_clock[2] ),
    .A3(\mod.div_clock[3] ),
    .S0(net27),
    .S1(net1),
    .X(_146_));
 sky130_fd_sc_hd__clkbuf_1 _264_ (.A(_146_),
    .X(\mod.clock_syn ));
 sky130_fd_sc_hd__inv_2 _265_ (.A(net7),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(net6),
    .Y(_148_));
 sky130_fd_sc_hd__o22a_1 _267_ (.A1(\mod.clock_counter_a[5] ),
    .A2(_147_),
    .B1(_148_),
    .B2(\mod.clock_counter_a[4] ),
    .X(_149_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(net4),
    .Y(_150_));
 sky130_fd_sc_hd__or2b_1 _269_ (.A(\mod.clock_counter_a[1] ),
    .B_N(net3),
    .X(_151_));
 sky130_fd_sc_hd__and2b_1 _270_ (.A_N(net2),
    .B(\mod.clock_counter_a[0] ),
    .X(_152_));
 sky130_fd_sc_hd__and2b_1 _271_ (.A_N(net3),
    .B(\mod.clock_counter_a[1] ),
    .X(_032_));
 sky130_fd_sc_hd__a221o_1 _272_ (.A1(\mod.clock_counter_a[2] ),
    .A2(_150_),
    .B1(_151_),
    .B2(_152_),
    .C1(_032_),
    .X(_033_));
 sky130_fd_sc_hd__inv_2 _273_ (.A(net5),
    .Y(_034_));
 sky130_fd_sc_hd__o22a_1 _274_ (.A1(\mod.clock_counter_a[3] ),
    .A2(_034_),
    .B1(_150_),
    .B2(\mod.clock_counter_a[2] ),
    .X(_035_));
 sky130_fd_sc_hd__a22o_1 _275_ (.A1(\mod.clock_counter_a[4] ),
    .A2(_148_),
    .B1(_034_),
    .B2(\mod.clock_counter_a[3] ),
    .X(_036_));
 sky130_fd_sc_hd__a21o_1 _276_ (.A1(_033_),
    .A2(_035_),
    .B1(_036_),
    .X(_037_));
 sky130_fd_sc_hd__a221oi_4 _277_ (.A1(\mod.clock_counter_a[5] ),
    .A2(_147_),
    .B1(_149_),
    .B2(_037_),
    .C1(\mod.clock_counter_a[6] ),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_1 _278_ (.A(\mod.div_clock[0] ),
    .B(_038_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(net13),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(net12),
    .Y(_040_));
 sky130_fd_sc_hd__o22a_1 _281_ (.A1(\mod.clock_counter_b[5] ),
    .A2(_039_),
    .B1(_040_),
    .B2(\mod.clock_counter_b[4] ),
    .X(_041_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(net10),
    .Y(_042_));
 sky130_fd_sc_hd__or2b_1 _283_ (.A(\mod.clock_counter_b[1] ),
    .B_N(net9),
    .X(_043_));
 sky130_fd_sc_hd__and2b_1 _284_ (.A_N(net8),
    .B(\mod.clock_counter_b[0] ),
    .X(_044_));
 sky130_fd_sc_hd__and2b_1 _285_ (.A_N(net9),
    .B(\mod.clock_counter_b[1] ),
    .X(_045_));
 sky130_fd_sc_hd__a221o_1 _286_ (.A1(\mod.clock_counter_b[2] ),
    .A2(_042_),
    .B1(_043_),
    .B2(_044_),
    .C1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(net11),
    .Y(_047_));
 sky130_fd_sc_hd__o22a_1 _288_ (.A1(\mod.clock_counter_b[3] ),
    .A2(_047_),
    .B1(_042_),
    .B2(\mod.clock_counter_b[2] ),
    .X(_048_));
 sky130_fd_sc_hd__a22o_1 _289_ (.A1(\mod.clock_counter_b[4] ),
    .A2(_040_),
    .B1(_047_),
    .B2(\mod.clock_counter_b[3] ),
    .X(_049_));
 sky130_fd_sc_hd__a21o_1 _290_ (.A1(_046_),
    .A2(_048_),
    .B1(_049_),
    .X(_050_));
 sky130_fd_sc_hd__a221oi_4 _291_ (.A1(\mod.clock_counter_b[5] ),
    .A2(_039_),
    .B1(_041_),
    .B2(_050_),
    .C1(\mod.clock_counter_b[6] ),
    .Y(_051_));
 sky130_fd_sc_hd__xnor2_1 _292_ (.A(\mod.div_clock[1] ),
    .B(_051_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(net19),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(net18),
    .Y(_053_));
 sky130_fd_sc_hd__o22a_1 _295_ (.A1(\mod.clock_counter_c[5] ),
    .A2(_052_),
    .B1(_053_),
    .B2(\mod.clock_counter_c[4] ),
    .X(_054_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(net16),
    .Y(_055_));
 sky130_fd_sc_hd__or2b_1 _297_ (.A(\mod.clock_counter_c[1] ),
    .B_N(net15),
    .X(_056_));
 sky130_fd_sc_hd__and2b_1 _298_ (.A_N(net14),
    .B(\mod.clock_counter_c[0] ),
    .X(_057_));
 sky130_fd_sc_hd__and2b_1 _299_ (.A_N(net15),
    .B(\mod.clock_counter_c[1] ),
    .X(_058_));
 sky130_fd_sc_hd__a221o_1 _300_ (.A1(\mod.clock_counter_c[2] ),
    .A2(_055_),
    .B1(_056_),
    .B2(_057_),
    .C1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(net17),
    .Y(_060_));
 sky130_fd_sc_hd__o22a_1 _302_ (.A1(\mod.clock_counter_c[3] ),
    .A2(_060_),
    .B1(_055_),
    .B2(\mod.clock_counter_c[2] ),
    .X(_061_));
 sky130_fd_sc_hd__a22o_1 _303_ (.A1(\mod.clock_counter_c[4] ),
    .A2(_053_),
    .B1(_060_),
    .B2(\mod.clock_counter_c[3] ),
    .X(_062_));
 sky130_fd_sc_hd__a21o_1 _304_ (.A1(_059_),
    .A2(_061_),
    .B1(_062_),
    .X(_063_));
 sky130_fd_sc_hd__a221oi_4 _305_ (.A1(\mod.clock_counter_c[5] ),
    .A2(_052_),
    .B1(_054_),
    .B2(_063_),
    .C1(\mod.clock_counter_c[6] ),
    .Y(_064_));
 sky130_fd_sc_hd__xnor2_1 _306_ (.A(\mod.div_clock[2] ),
    .B(_064_),
    .Y(_002_));
 sky130_fd_sc_hd__dfxtp_1 _307_ (.CLK(net32),
    .D(_000_),
    .Q(\mod.div_clock[0] ));
 sky130_fd_sc_hd__dfxtp_1 _308_ (.CLK(net30),
    .D(_001_),
    .Q(\mod.div_clock[1] ));
 sky130_fd_sc_hd__dfxtp_1 _309_ (.CLK(net30),
    .D(_002_),
    .Q(\mod.div_clock[2] ));
 sky130_fd_sc_hd__dfxtp_1 _310_ (.CLK(net30),
    .D(_003_),
    .Q(\mod.div_clock[3] ));
 sky130_fd_sc_hd__dfxtp_1 _311_ (.CLK(net29),
    .D(_004_),
    .Q(\mod.clock_counter_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _312_ (.CLK(net29),
    .D(_005_),
    .Q(\mod.clock_counter_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _313_ (.CLK(net29),
    .D(_006_),
    .Q(\mod.clock_counter_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _314_ (.CLK(net29),
    .D(_007_),
    .Q(\mod.clock_counter_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _315_ (.CLK(net29),
    .D(_008_),
    .Q(\mod.clock_counter_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _316_ (.CLK(net29),
    .D(_009_),
    .Q(\mod.clock_counter_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _317_ (.CLK(net29),
    .D(_010_),
    .Q(\mod.clock_counter_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _318_ (.CLK(net29),
    .D(_011_),
    .Q(\mod.clock_counter_c[0] ));
 sky130_fd_sc_hd__dfxtp_1 _319_ (.CLK(net29),
    .D(_012_),
    .Q(\mod.clock_counter_c[1] ));
 sky130_fd_sc_hd__dfxtp_1 _320_ (.CLK(net29),
    .D(_013_),
    .Q(\mod.clock_counter_c[2] ));
 sky130_fd_sc_hd__dfxtp_1 _321_ (.CLK(net30),
    .D(_014_),
    .Q(\mod.clock_counter_c[3] ));
 sky130_fd_sc_hd__dfxtp_1 _322_ (.CLK(net30),
    .D(_015_),
    .Q(\mod.clock_counter_c[4] ));
 sky130_fd_sc_hd__dfxtp_1 _323_ (.CLK(net30),
    .D(_016_),
    .Q(\mod.clock_counter_c[5] ));
 sky130_fd_sc_hd__dfxtp_1 _324_ (.CLK(net30),
    .D(_017_),
    .Q(\mod.clock_counter_c[6] ));
 sky130_fd_sc_hd__dfxtp_1 _325_ (.CLK(net30),
    .D(_018_),
    .Q(\mod.clock_counter_b[0] ));
 sky130_fd_sc_hd__dfxtp_1 _326_ (.CLK(net30),
    .D(_019_),
    .Q(\mod.clock_counter_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _327_ (.CLK(net31),
    .D(_020_),
    .Q(\mod.clock_counter_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _328_ (.CLK(net31),
    .D(_021_),
    .Q(\mod.clock_counter_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _329_ (.CLK(net31),
    .D(_022_),
    .Q(\mod.clock_counter_b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _330_ (.CLK(net31),
    .D(_023_),
    .Q(\mod.clock_counter_b[5] ));
 sky130_fd_sc_hd__dfxtp_1 _331_ (.CLK(net31),
    .D(_024_),
    .Q(\mod.clock_counter_b[6] ));
 sky130_fd_sc_hd__dfxtp_1 _332_ (.CLK(net32),
    .D(_025_),
    .Q(\mod.clock_counter_a[0] ));
 sky130_fd_sc_hd__dfxtp_1 _333_ (.CLK(net32),
    .D(_026_),
    .Q(\mod.clock_counter_a[1] ));
 sky130_fd_sc_hd__dfxtp_1 _334_ (.CLK(net32),
    .D(_027_),
    .Q(\mod.clock_counter_a[2] ));
 sky130_fd_sc_hd__dfxtp_1 _335_ (.CLK(net32),
    .D(_028_),
    .Q(\mod.clock_counter_a[3] ));
 sky130_fd_sc_hd__dfxtp_1 _336_ (.CLK(net32),
    .D(_029_),
    .Q(\mod.clock_counter_a[4] ));
 sky130_fd_sc_hd__dfxtp_1 _337_ (.CLK(net32),
    .D(_030_),
    .Q(\mod.clock_counter_a[5] ));
 sky130_fd_sc_hd__dfxtp_1 _338_ (.CLK(net32),
    .D(_031_),
    .Q(\mod.clock_counter_a[6] ));
 sky130_fd_sc_hd__conb_1 tiny_user_project_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tiny_user_project_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tiny_user_project_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tiny_user_project_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tiny_user_project_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tiny_user_project_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tiny_user_project_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tiny_user_project_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tiny_user_project_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tiny_user_project_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tiny_user_project_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tiny_user_project_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 tiny_user_project_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 tiny_user_project_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 tiny_user_project_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tiny_user_project_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tiny_user_project_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tiny_user_project_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tiny_user_project_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tiny_user_project_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tiny_user_project_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tiny_user_project_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tiny_user_project_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tiny_user_project_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tiny_user_project_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tiny_user_project_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tiny_user_project_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tiny_user_project_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tiny_user_project_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tiny_user_project_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tiny_user_project_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tiny_user_project_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tiny_user_project_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tiny_user_project_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tiny_user_project_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tiny_user_project_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tiny_user_project_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tiny_user_project_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tiny_user_project_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tiny_user_project_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tiny_user_project_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tiny_user_project_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tiny_user_project_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tiny_user_project_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 tiny_user_project_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 tiny_user_project_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 tiny_user_project_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 tiny_user_project_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 tiny_user_project_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 tiny_user_project_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 tiny_user_project_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 tiny_user_project_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 tiny_user_project_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 tiny_user_project_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 tiny_user_project_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 tiny_user_project_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 tiny_user_project_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 tiny_user_project_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 tiny_user_project_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 tiny_user_project_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 tiny_user_project_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 tiny_user_project_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 tiny_user_project_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 tiny_user_project_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 tiny_user_project_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 tiny_user_project_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 tiny_user_project_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 tiny_user_project_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 tiny_user_project_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 tiny_user_project_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 tiny_user_project_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 tiny_user_project_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 tiny_user_project_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 tiny_user_project_107 (.LO(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[10]));
 sky130_fd_sc_hd__clkbuf_1 _414_ (.A(\mod.clock_syn ),
    .X(net28));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[10]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[11]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[12]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[13]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[14]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[16]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(io_in[17]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(io_in[18]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[19]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[20]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(io_in[21]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[22]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(io_in[23]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(io_in[24]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(io_in[25]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(io_in[26]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(io_in[27]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(io_in[28]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(io_in[29]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(io_in[30]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(io_in[31]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(io_in[32]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(io_in[33]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(io_in[34]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(io_in[8]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(io_in[9]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[35]));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net26),
    .X(net32));
 sky130_fd_sc_hd__conb_1 tiny_user_project_33 (.LO(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_188 ();
 assign io_oeb[0] = net33;
 assign io_oeb[10] = net43;
 assign io_oeb[11] = net44;
 assign io_oeb[12] = net45;
 assign io_oeb[13] = net46;
 assign io_oeb[14] = net47;
 assign io_oeb[15] = net48;
 assign io_oeb[16] = net49;
 assign io_oeb[17] = net50;
 assign io_oeb[18] = net51;
 assign io_oeb[19] = net52;
 assign io_oeb[1] = net34;
 assign io_oeb[20] = net53;
 assign io_oeb[21] = net54;
 assign io_oeb[22] = net55;
 assign io_oeb[23] = net56;
 assign io_oeb[24] = net57;
 assign io_oeb[25] = net58;
 assign io_oeb[26] = net59;
 assign io_oeb[27] = net60;
 assign io_oeb[28] = net61;
 assign io_oeb[29] = net62;
 assign io_oeb[2] = net35;
 assign io_oeb[30] = net63;
 assign io_oeb[31] = net64;
 assign io_oeb[32] = net65;
 assign io_oeb[33] = net66;
 assign io_oeb[34] = net67;
 assign io_oeb[35] = net68;
 assign io_oeb[36] = net69;
 assign io_oeb[37] = net70;
 assign io_oeb[3] = net36;
 assign io_oeb[4] = net37;
 assign io_oeb[5] = net38;
 assign io_oeb[6] = net39;
 assign io_oeb[7] = net40;
 assign io_oeb[8] = net41;
 assign io_oeb[9] = net42;
 assign io_out[0] = net71;
 assign io_out[10] = net81;
 assign io_out[11] = net82;
 assign io_out[12] = net83;
 assign io_out[13] = net84;
 assign io_out[14] = net85;
 assign io_out[15] = net86;
 assign io_out[16] = net87;
 assign io_out[17] = net88;
 assign io_out[18] = net89;
 assign io_out[19] = net90;
 assign io_out[1] = net72;
 assign io_out[20] = net91;
 assign io_out[21] = net92;
 assign io_out[22] = net93;
 assign io_out[23] = net94;
 assign io_out[24] = net95;
 assign io_out[25] = net96;
 assign io_out[26] = net97;
 assign io_out[27] = net98;
 assign io_out[28] = net99;
 assign io_out[29] = net100;
 assign io_out[2] = net73;
 assign io_out[30] = net101;
 assign io_out[31] = net102;
 assign io_out[32] = net103;
 assign io_out[33] = net104;
 assign io_out[34] = net105;
 assign io_out[36] = net106;
 assign io_out[37] = net107;
 assign io_out[3] = net74;
 assign io_out[4] = net75;
 assign io_out[5] = net76;
 assign io_out[6] = net77;
 assign io_out[7] = net78;
 assign io_out[8] = net79;
 assign io_out[9] = net80;
endmodule

